`timescale 1 ns / 1 ns module xRgm1KQSpBEMURvTRAnYsB (v04pHKxyc2sPW047bbyUgE, JAMOfrNHxGSYDF0urqkLN, Ebx0yJLDGKevxkqzRPIfvG, B58twvtfgVWGK5P29KavtH, qhk6Uhwhppvpssqm7Nh6XE, VWSiqDgxQN9a2J7zRy3p4E, LhqlKpPzANkuN2xC8HYciC, jNZ4xylBKAANfCL11XNxzB, R6zf5iqRNVEGVBO8egq8kF, A5SQIaNgqW7DcTqQkKRVeD, GaetbCaMty7UkzjqNoYErC, k3VfrgkD6DWITJL9WW5W4D, pPn6MVGqBLqJ0xzN2WYfFG, Pq4nKEqqr18aLXK1kX1dfH); input v04pHKxyc2sPW047bbyUgE; input JAMOfrNHxGSYDF0urqkLN; input Ebx0yJLDGKevxkqzRPIfvG; input signed [15:0] B58twvtfgVWGK5P29KavtH; input signed [15:0] qhk6Uhwhppvpssqm7Nh6XE; input signed [15:0] VWSiqDgxQN9a2J7zRy3p4E; input signed [15:0] LhqlKpPzANkuN2xC8HYciC; input jNZ4xylBKAANfCL11XNxzB; input R6zf5iqRNVEGVBO8egq8kF; output signed [15:0] A5SQIaNgqW7DcTqQkKRVeD; output signed [15:0] GaetbCaMty7UkzjqNoYErC; output signed [15:0] k3VfrgkD6DWITJL9WW5W4D; output signed [15:0] pPn6MVGqBLqJ0xzN2WYfFG; output Pq4nKEqqr18aLXK1kX1dfH; reg AxdzJminNkFCybtxxeC5hH; reg signed [16:0] p9Q1ZdD8IyrQGhwT1XXpAwH; reg signed [16:0] FrouE4YVttOqChzztq9MRG; reg signed [16:0] i4FJCC6Xft9yUijVwpyTC0E; reg signed [16:0] N5RqGyuQKrj2dkBK5NIpfD; reg b8PGIsG3FsdAJqb7hOUD1oC; reg signed [16:0] u6qmTF9ijEkH9xmDrm95pEF; reg signed [16:0] MP4qvH0uMShcprYVFxKkUD; reg signed [16:0] COyf11G22yt2ahr9Ucug2E; reg signed [16:0] bYOlGODgGA4hK2uJ9g4xaG; reg signed [15:0] wzDrz6Bb4WkvBDnpgbSZ9E; reg signed [15:0] rddvPMIplivXE2pWkXTaQB; reg signed [15:0] M5AqS9R7rFTkWxwo8io2rH; reg signed [15:0] lcJo4MnEaj41ofRAtLkn4D; reg z4CQk9lB9oVzTWAolXGwv3G; reg signed [16:0] a6WUK3shR7OoXJD6OQBcnbC; reg signed [16:0] z8sdLNMywEyzxM9eSpPklMB; reg signed [16:0] x4JZ8sOjxjZWNeN08B95t5B; reg signed [16:0] JpNj7HaVF5ISgAz8d6xCmE; reg signed [16:0] lyJA6GgUdA5yMT3KGmkiBB; reg signed [16:0] YTn6r1K2cbi4BzelKHgZMH; reg signed [16:0] T6fhnGgnCx4gzNMLRlfJsB; reg signed [16:0] QaUWOROgNo7uvlOzzIL7gF; reg signed [16:0] f9uiVizQ8iG3TggFQMEaqMB; reg signed [16:0] whyOPXTaiRJEg5hgsaLJCG; reg signed [16:0] yqGXdE6pHXRFGlXkfvbpKC; reg signed [16:0] UzOnWFVNmsGSUzlrKfHqwF; reg signed [16:0] b9p1O84anZ1REVMvdH9T6cE; reg signed [16:0] uOyZcxygSH2ObqTFvmjZLD; reg signed [16:0] giifcHhQs1eZ2W9VasanfG; reg signed [16:0] Ht14IixEv7IQddUNB8FBaF; reg signed [16:0] g64FBA6XTYfJB3gQdH04OJH; reg signed [16:0] cefQ41MlYs7FI4dPMnads; reg signed [16:0] ZLjCoy1mhX7nS8r36AkTnG; reg signed [16:0] z6qazKI7KMGAFLe2KGVVFE; reg signed [16:0] xE4ft4QLMQrp1NtpcdoU2D; reg signed [16:0] b3b6q6yOnUzkdBZha4J35NB; reg signed [16:0] xsDfZ2jarysSjALlotRtW; reg signed [16:0] YLWHYhSBwDrFHhQzmw106G; reg signed [16:0] J3I5o2R6c9ixHmw1Oa9EvE; reg signed [16:0] bN7pv94LbbUjIRAxJt4lf; reg signed [16:0] PZRWIojv1r4p0mRa5bnL8G; reg signed [16:0] iZxjhcD6M6J4jJWVBLDvjG; wire al5EhrIEQ1yUUqlDvo19NC; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : aMdxH72OgWBZw20gQc6DxE if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin AxdzJminNkFCybtxxeC5hH <= 1'b0; p9Q1ZdD8IyrQGhwT1XXpAwH <= 17'sb00000000000000000; FrouE4YVttOqChzztq9MRG <= 17'sb00000000000000000; i4FJCC6Xft9yUijVwpyTC0E <= 17'sb00000000000000000; N5RqGyuQKrj2dkBK5NIpfD <= 17'sb00000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin AxdzJminNkFCybtxxeC5hH <= 1'b0; p9Q1ZdD8IyrQGhwT1XXpAwH <= 17'sb00000000000000000; FrouE4YVttOqChzztq9MRG <= 17'sb00000000000000000; i4FJCC6Xft9yUijVwpyTC0E <= 17'sb00000000000000000; N5RqGyuQKrj2dkBK5NIpfD <= 17'sb00000000000000000; end else begin AxdzJminNkFCybtxxeC5hH <= b8PGIsG3FsdAJqb7hOUD1oC; p9Q1ZdD8IyrQGhwT1XXpAwH <= u6qmTF9ijEkH9xmDrm95pEF; FrouE4YVttOqChzztq9MRG <= MP4qvH0uMShcprYVFxKkUD; i4FJCC6Xft9yUijVwpyTC0E <= COyf11G22yt2ahr9Ucug2E; N5RqGyuQKrj2dkBK5NIpfD <= bYOlGODgGA4hK2uJ9g4xaG; end end end always @(AxdzJminNkFCybtxxeC5hH, B58twvtfgVWGK5P29KavtH, Ebx0yJLDGKevxkqzRPIfvG, FrouE4YVttOqChzztq9MRG, LhqlKpPzANkuN2xC8HYciC, N5RqGyuQKrj2dkBK5NIpfD, VWSiqDgxQN9a2J7zRy3p4E, i4FJCC6Xft9yUijVwpyTC0E, jNZ4xylBKAANfCL11XNxzB, p9Q1ZdD8IyrQGhwT1XXpAwH, qhk6Uhwhppvpssqm7Nh6XE) begin b9p1O84anZ1REVMvdH9T6cE = 17'sb00000000000000000; uOyZcxygSH2ObqTFvmjZLD = 17'sb00000000000000000; giifcHhQs1eZ2W9VasanfG = 17'sb00000000000000000; Ht14IixEv7IQddUNB8FBaF = 17'sb00000000000000000; g64FBA6XTYfJB3gQdH04OJH = 17'sb00000000000000000; cefQ41MlYs7FI4dPMnads = 17'sb00000000000000000; ZLjCoy1mhX7nS8r36AkTnG = 17'sb00000000000000000; z6qazKI7KMGAFLe2KGVVFE = 17'sb00000000000000000; xE4ft4QLMQrp1NtpcdoU2D = 17'sb00000000000000000; b3b6q6yOnUzkdBZha4J35NB = 17'sb00000000000000000; xsDfZ2jarysSjALlotRtW = 17'sb00000000000000000; YLWHYhSBwDrFHhQzmw106G = 17'sb00000000000000000; J3I5o2R6c9ixHmw1Oa9EvE = 17'sb00000000000000000; bN7pv94LbbUjIRAxJt4lf = 17'sb00000000000000000; PZRWIojv1r4p0mRa5bnL8G = 17'sb00000000000000000; iZxjhcD6M6J4jJWVBLDvjG = 17'sb00000000000000000; u6qmTF9ijEkH9xmDrm95pEF = p9Q1ZdD8IyrQGhwT1XXpAwH; MP4qvH0uMShcprYVFxKkUD = FrouE4YVttOqChzztq9MRG; COyf11G22yt2ahr9Ucug2E = i4FJCC6Xft9yUijVwpyTC0E; bYOlGODgGA4hK2uJ9g4xaG = N5RqGyuQKrj2dkBK5NIpfD; b8PGIsG3FsdAJqb7hOUD1oC = jNZ4xylBKAANfCL11XNxzB; if (Ebx0yJLDGKevxkqzRPIfvG != 1'b0) begin if (jNZ4xylBKAANfCL11XNxzB) begin b9p1O84anZ1REVMvdH9T6cE = {B58twvtfgVWGK5P29KavtH[15], B58twvtfgVWGK5P29KavtH}; uOyZcxygSH2ObqTFvmjZLD = {LhqlKpPzANkuN2xC8HYciC[15], LhqlKpPzANkuN2xC8HYciC}; u6qmTF9ijEkH9xmDrm95pEF = b9p1O84anZ1REVMvdH9T6cE + uOyZcxygSH2ObqTFvmjZLD; giifcHhQs1eZ2W9VasanfG = {B58twvtfgVWGK5P29KavtH[15], B58twvtfgVWGK5P29KavtH}; Ht14IixEv7IQddUNB8FBaF = {LhqlKpPzANkuN2xC8HYciC[15], LhqlKpPzANkuN2xC8HYciC}; COyf11G22yt2ahr9Ucug2E = giifcHhQs1eZ2W9VasanfG - Ht14IixEv7IQddUNB8FBaF; g64FBA6XTYfJB3gQdH04OJH = {qhk6Uhwhppvpssqm7Nh6XE[15], qhk6Uhwhppvpssqm7Nh6XE}; cefQ41MlYs7FI4dPMnads = {VWSiqDgxQN9a2J7zRy3p4E[15], VWSiqDgxQN9a2J7zRy3p4E}; bYOlGODgGA4hK2uJ9g4xaG = g64FBA6XTYfJB3gQdH04OJH + cefQ41MlYs7FI4dPMnads; ZLjCoy1mhX7nS8r36AkTnG = {qhk6Uhwhppvpssqm7Nh6XE[15], qhk6Uhwhppvpssqm7Nh6XE}; z6qazKI7KMGAFLe2KGVVFE = {VWSiqDgxQN9a2J7zRy3p4E[15], VWSiqDgxQN9a2J7zRy3p4E}; MP4qvH0uMShcprYVFxKkUD = ZLjCoy1mhX7nS8r36AkTnG - z6qazKI7KMGAFLe2KGVVFE; end end else if (jNZ4xylBKAANfCL11XNxzB) begin xE4ft4QLMQrp1NtpcdoU2D = {B58twvtfgVWGK5P29KavtH[15], B58twvtfgVWGK5P29KavtH}; b3b6q6yOnUzkdBZha4J35NB = {VWSiqDgxQN9a2J7zRy3p4E[15], VWSiqDgxQN9a2J7zRy3p4E}; u6qmTF9ijEkH9xmDrm95pEF = xE4ft4QLMQrp1NtpcdoU2D + b3b6q6yOnUzkdBZha4J35NB; xsDfZ2jarysSjALlotRtW = {B58twvtfgVWGK5P29KavtH[15], B58twvtfgVWGK5P29KavtH}; YLWHYhSBwDrFHhQzmw106G = {VWSiqDgxQN9a2J7zRy3p4E[15], VWSiqDgxQN9a2J7zRy3p4E}; COyf11G22yt2ahr9Ucug2E = xsDfZ2jarysSjALlotRtW - YLWHYhSBwDrFHhQzmw106G; J3I5o2R6c9ixHmw1Oa9EvE = {qhk6Uhwhppvpssqm7Nh6XE[15], qhk6Uhwhppvpssqm7Nh6XE}; bN7pv94LbbUjIRAxJt4lf = {LhqlKpPzANkuN2xC8HYciC[15], LhqlKpPzANkuN2xC8HYciC}; MP4qvH0uMShcprYVFxKkUD = J3I5o2R6c9ixHmw1Oa9EvE + bN7pv94LbbUjIRAxJt4lf; PZRWIojv1r4p0mRa5bnL8G = {qhk6Uhwhppvpssqm7Nh6XE[15], qhk6Uhwhppvpssqm7Nh6XE}; iZxjhcD6M6J4jJWVBLDvjG = {LhqlKpPzANkuN2xC8HYciC[15], LhqlKpPzANkuN2xC8HYciC}; bYOlGODgGA4hK2uJ9g4xaG = PZRWIojv1r4p0mRa5bnL8G - iZxjhcD6M6J4jJWVBLDvjG; end a6WUK3shR7OoXJD6OQBcnbC = ({p9Q1ZdD8IyrQGhwT1XXpAwH[16], p9Q1ZdD8IyrQGhwT1XXpAwH[16:1]}) + $signed({1'b0, p9Q1ZdD8IyrQGhwT1XXpAwH[0]}); z8sdLNMywEyzxM9eSpPklMB = a6WUK3shR7OoXJD6OQBcnbC >>> 8'd1; x4JZ8sOjxjZWNeN08B95t5B = {z8sdLNMywEyzxM9eSpPklMB[15:0], 1'b0}; wzDrz6Bb4WkvBDnpgbSZ9E = x4JZ8sOjxjZWNeN08B95t5B[15:0]; JpNj7HaVF5ISgAz8d6xCmE = ({FrouE4YVttOqChzztq9MRG[16], FrouE4YVttOqChzztq9MRG[16:1]}) + $signed({1'b0, FrouE4YVttOqChzztq9MRG[0]}); lyJA6GgUdA5yMT3KGmkiBB = JpNj7HaVF5ISgAz8d6xCmE >>> 8'd1; YTn6r1K2cbi4BzelKHgZMH = {lyJA6GgUdA5yMT3KGmkiBB[15:0], 1'b0}; rddvPMIplivXE2pWkXTaQB = YTn6r1K2cbi4BzelKHgZMH[15:0]; T6fhnGgnCx4gzNMLRlfJsB = ({i4FJCC6Xft9yUijVwpyTC0E[16], i4FJCC6Xft9yUijVwpyTC0E[16:1]}) + $signed({1'b0, i4FJCC6Xft9yUijVwpyTC0E[0]}); QaUWOROgNo7uvlOzzIL7gF = T6fhnGgnCx4gzNMLRlfJsB >>> 8'd1; f9uiVizQ8iG3TggFQMEaqMB = {QaUWOROgNo7uvlOzzIL7gF[15:0], 1'b0}; M5AqS9R7rFTkWxwo8io2rH = f9uiVizQ8iG3TggFQMEaqMB[15:0]; whyOPXTaiRJEg5hgsaLJCG = ({N5RqGyuQKrj2dkBK5NIpfD[16], N5RqGyuQKrj2dkBK5NIpfD[16:1]}) + $signed({1'b0, N5RqGyuQKrj2dkBK5NIpfD[0]}); yqGXdE6pHXRFGlXkfvbpKC = whyOPXTaiRJEg5hgsaLJCG >>> 8'd1; UzOnWFVNmsGSUzlrKfHqwF = {yqGXdE6pHXRFGlXkfvbpKC[15:0], 1'b0}; lcJo4MnEaj41ofRAtLkn4D = UzOnWFVNmsGSUzlrKfHqwF[15:0]; z4CQk9lB9oVzTWAolXGwv3G = AxdzJminNkFCybtxxeC5hH; end assign A5SQIaNgqW7DcTqQkKRVeD = wzDrz6Bb4WkvBDnpgbSZ9E; assign GaetbCaMty7UkzjqNoYErC = rddvPMIplivXE2pWkXTaQB; assign k3VfrgkD6DWITJL9WW5W4D = M5AqS9R7rFTkWxwo8io2rH; assign pPn6MVGqBLqJ0xzN2WYfFG = lcJo4MnEaj41ofRAtLkn4D; assign Pq4nKEqqr18aLXK1kX1dfH = z4CQk9lB9oVzTWAolXGwv3G; endmodule