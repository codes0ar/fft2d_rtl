`timescale 1 ns / 1 ns module xhnyoB96GyFxIQr6c1oc4G (v04pHKxyc2sPW047bbyUgE, JAMOfrNHxGSYDF0urqkLN, JdpDaA8gpSp0rE35OGZkGE, mgknRxAcgFrHqTt5CZvnSF, sCFM4WicR6deeSAdSwumP, BKNY6GzA6oGZumjzTATycD, uUcj3UAzjmPW47yNyzbT8C, uwZv0qzQLi0MDBWLWzKuAG, n65LdbEr6NMNaEFcjX8Fh6F, x9j7a5gok64zzNKnvdJNnE, bPL0FcLvoxhO0amTUOV9QC, r4JngA0ZVhEElGRZci9fohF, a8xx20Fc5nKc8DbqSwNBuB, vLT6ef7BJliTDpt4k5jqF, R6zf5iqRNVEGVBO8egq8kF, N2ZdE4zLlq5uRV4rcE2wdE, AECH0r3KnKo0RJFepDhYUD, twcuYIJzeZMBjyHmZ1FZDD, f3NrgRvCkMfwf1E3PnKtczF, f2XZKbXdctKWPTTQYeLkBWE); input v04pHKxyc2sPW047bbyUgE; input JAMOfrNHxGSYDF0urqkLN; input JdpDaA8gpSp0rE35OGZkGE; input signed [15:0] mgknRxAcgFrHqTt5CZvnSF; input signed [15:0] sCFM4WicR6deeSAdSwumP; input BKNY6GzA6oGZumjzTATycD; input signed [15:0] uUcj3UAzjmPW47yNyzbT8C; input signed [15:0] uwZv0qzQLi0MDBWLWzKuAG; input n65LdbEr6NMNaEFcjX8Fh6F; input signed [15:0] x9j7a5gok64zzNKnvdJNnE; input signed [15:0] bPL0FcLvoxhO0amTUOV9QC; input signed [15:0] r4JngA0ZVhEElGRZci9fohF; input signed [15:0] a8xx20Fc5nKc8DbqSwNBuB; input vLT6ef7BJliTDpt4k5jqF; input R6zf5iqRNVEGVBO8egq8kF; output signed [15:0] N2ZdE4zLlq5uRV4rcE2wdE; output [6:0] AECH0r3KnKo0RJFepDhYUD; output twcuYIJzeZMBjyHmZ1FZDD; output signed [15:0] f3NrgRvCkMfwf1E3PnKtczF; output signed [15:0] f2XZKbXdctKWPTTQYeLkBWE; reg signed [15:0] ERpxhnx4yQO2gF4g0J9G8G; reg signed [15:0] yAfJq6fAufU3HOal8Q4DkG; reg yeHXFGHVMgEtZ4f1O7U2OB; reg [6:0] w7JAMsElgYTLo8syEMZ8Lk; reg [2:0] skXEjqLZnGZAr6RJ8QjjD; reg [1:0] r2jaHd7wMNX07DmqtoTGYfB; reg [6:0] MDWW9wjzQsTkpJTsAXw1tG; reg signed [15:0] CDiyyho6hDs0nvcIRHvdfF; reg signed [15:0] EIQhCDitCjjxqIfp1PqavH; reg PRVmCVU2hynJRxCDsjx8OE; reg signed [15:0] l96dMLSJZGbzKOOaSawmDC; reg signed [15:0] h7QHiA6jfRB0V5iS7nYrsR; reg [2:0] pN9XTk8HB1jtfigsDxuKfE; reg ucLx3e73qDSgpZETH1oJ9; reg [2:0] BAQ1YrOPn1tEt43kT1QPvE; reg [2:0] oFHbC0LQKaxvW8gPAQzBAB; reg yUuRVFmKCNYKHMIon8qCKG; reg c1qRGYMEWodUPO7ZFq831QB; reg OTCxoIqhEhA65VRuJvFoxB; reg signed [15:0] U2JXBqjMcwW1AxVU5Q1ESG; reg signed [15:0] bm6UZNfjlfNI5cDV8oaTj; reg EzzigQlTGv8J7DBTRmqQ9C; reg [6:0] srDEOQxwGboahrxQGs2vYE; reg [2:0] gZNZkxioohAMHXxms1BEOE; reg [1:0] xhZyruBklMjVnVQHFCsnC; reg [6:0] MTuGLzs6sZnejyrpSaOMvF; reg signed [15:0] tArVqL2CTwuHoaoeSuZkaB; reg signed [15:0] g4P4JTWbBBBn0JhReP8eXAH; reg f1bIHzdG7kDHnL70sxnVWzB; reg signed [15:0] s3m9T9rV2e4ZoMyZFS4lKeB; reg signed [15:0] p7ixx7ZWknoF1F7FbI5yjED; reg [2:0] KwC6wbRFLWpjZZERCcYIGB; reg MOh79n10Ewq3O8I6VYlcS; reg [2:0] Ym7Bnv0nBa8mPH5deUne6F; reg [2:0] e2MNnweVMUgzBGV1fQxq5dB; reg A9eIucMmprrI3z0XPuKfq; reg CdyHxmDTkJd4Kce0MGL8uE; reg BlSFAnc8BhBCmuAIbP8voB; reg signed [15:0] r5kivPzvWgOSiA0gZBDsCMD; reg signed [15:0] iOhy3XYM3su7ndksftfCZG; reg [6:0] TIIVgGzxbljXJKElx1RmZB; reg d4GqKaFZXLUlts9HBCZPXG; reg signed [15:0] lJc3nzBSuIub4Fgm41LhsH; reg signed [15:0] e4s7lktq7sxpTrarrx3LfPD; reg [2:0] mmaX8nGKzNYVdRyx6p1LtC; reg whMUFL1J2R7VsHTN9UxHOH; reg [2:0] pfAgd4CSuF40Tz4AXQRjjB; reg tKu1I9axj5Jgdz0Uq0pTPF; reg signed [15:0] rM5MTP4UKZC3il6lMwiHT; reg signed [15:0] gP6GlHEmSHKO19LfKcs3AH; reg wyxMTJhenZ0YDgDbHfiMlC; wire signed [15:0] PLGAQRVd1M1QgFrsMrWVBH; wire signed [15:0] LifjwIUema6BHVuDJV77JF; reg signed [15:0] cWUwraq7WjwtV5SP0dQobH; reg signed [15:0] v1iHIP96KWtHSOQsfIP0oDD; reg r1RjufPwJY8CeBEsvwJ2flF; reg signed [15:0] HVkI4mR4uVjbZBmf8GvOyF; reg signed [15:0] VZmPcFtZLayUEhrt70JPkG; reg o59gL1lKXL2dKgQPA064uXG; reg signed [15:0] P3F2cuYaLRQxlfxwGBfSjF; reg signed [15:0] Rwrw0YN1HJLlhEzt1YbmaC; reg vl2rwYFSlP59iBJIjf8F4D; wire WYGJe9qM2amuIe1VNiR9e; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : N7A9w81SChJNEuxavvBOiF if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin ERpxhnx4yQO2gF4g0J9G8G <= 16'sb0000000000000000; yAfJq6fAufU3HOal8Q4DkG <= 16'sb0000000000000000; CDiyyho6hDs0nvcIRHvdfF <= 16'sb0000000000000000; EIQhCDitCjjxqIfp1PqavH <= 16'sb0000000000000000; PRVmCVU2hynJRxCDsjx8OE <= 1'b0; yeHXFGHVMgEtZ4f1O7U2OB <= 1'b0; skXEjqLZnGZAr6RJ8QjjD <= 3'b000; r2jaHd7wMNX07DmqtoTGYfB <= 2'b00; w7JAMsElgYTLo8syEMZ8Lk <= 7'b0000000; MDWW9wjzQsTkpJTsAXw1tG <= 7'b0000000; l96dMLSJZGbzKOOaSawmDC <= 16'sb0000000000000000; h7QHiA6jfRB0V5iS7nYrsR <= 16'sb0000000000000000; pN9XTk8HB1jtfigsDxuKfE <= 3'b000; ucLx3e73qDSgpZETH1oJ9 <= 1'b0; BAQ1YrOPn1tEt43kT1QPvE <= 3'b000; oFHbC0LQKaxvW8gPAQzBAB <= 3'b000; yUuRVFmKCNYKHMIon8qCKG <= 1'b0; c1qRGYMEWodUPO7ZFq831QB <= 1'b0; OTCxoIqhEhA65VRuJvFoxB <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin ERpxhnx4yQO2gF4g0J9G8G <= 16'sb0000000000000000; yAfJq6fAufU3HOal8Q4DkG <= 16'sb0000000000000000; CDiyyho6hDs0nvcIRHvdfF <= 16'sb0000000000000000; EIQhCDitCjjxqIfp1PqavH <= 16'sb0000000000000000; PRVmCVU2hynJRxCDsjx8OE <= 1'b0; yeHXFGHVMgEtZ4f1O7U2OB <= 1'b0; skXEjqLZnGZAr6RJ8QjjD <= 3'b000; r2jaHd7wMNX07DmqtoTGYfB <= 2'b00; w7JAMsElgYTLo8syEMZ8Lk <= 7'b0000000; MDWW9wjzQsTkpJTsAXw1tG <= 7'b0000000; l96dMLSJZGbzKOOaSawmDC <= 16'sb0000000000000000; h7QHiA6jfRB0V5iS7nYrsR <= 16'sb0000000000000000; pN9XTk8HB1jtfigsDxuKfE <= 3'b000; ucLx3e73qDSgpZETH1oJ9 <= 1'b0; BAQ1YrOPn1tEt43kT1QPvE <= 3'b000; oFHbC0LQKaxvW8gPAQzBAB <= 3'b000; yUuRVFmKCNYKHMIon8qCKG <= 1'b0; c1qRGYMEWodUPO7ZFq831QB <= 1'b0; OTCxoIqhEhA65VRuJvFoxB <= 1'b0; end else begin ERpxhnx4yQO2gF4g0J9G8G <= U2JXBqjMcwW1AxVU5Q1ESG; yAfJq6fAufU3HOal8Q4DkG <= bm6UZNfjlfNI5cDV8oaTj; yeHXFGHVMgEtZ4f1O7U2OB <= EzzigQlTGv8J7DBTRmqQ9C; w7JAMsElgYTLo8syEMZ8Lk <= srDEOQxwGboahrxQGs2vYE; skXEjqLZnGZAr6RJ8QjjD <= gZNZkxioohAMHXxms1BEOE; r2jaHd7wMNX07DmqtoTGYfB <= xhZyruBklMjVnVQHFCsnC; MDWW9wjzQsTkpJTsAXw1tG <= MTuGLzs6sZnejyrpSaOMvF; CDiyyho6hDs0nvcIRHvdfF <= tArVqL2CTwuHoaoeSuZkaB; EIQhCDitCjjxqIfp1PqavH <= g4P4JTWbBBBn0JhReP8eXAH; PRVmCVU2hynJRxCDsjx8OE <= f1bIHzdG7kDHnL70sxnVWzB; l96dMLSJZGbzKOOaSawmDC <= s3m9T9rV2e4ZoMyZFS4lKeB; h7QHiA6jfRB0V5iS7nYrsR <= p7ixx7ZWknoF1F7FbI5yjED; pN9XTk8HB1jtfigsDxuKfE <= KwC6wbRFLWpjZZERCcYIGB; ucLx3e73qDSgpZETH1oJ9 <= MOh79n10Ewq3O8I6VYlcS; BAQ1YrOPn1tEt43kT1QPvE <= Ym7Bnv0nBa8mPH5deUne6F; oFHbC0LQKaxvW8gPAQzBAB <= e2MNnweVMUgzBGV1fQxq5dB; yUuRVFmKCNYKHMIon8qCKG <= A9eIucMmprrI3z0XPuKfq; c1qRGYMEWodUPO7ZFq831QB <= CdyHxmDTkJd4Kce0MGL8uE; OTCxoIqhEhA65VRuJvFoxB <= BlSFAnc8BhBCmuAIbP8voB; end end end always @(BAQ1YrOPn1tEt43kT1QPvE, BKNY6GzA6oGZumjzTATycD, CDiyyho6hDs0nvcIRHvdfF, EIQhCDitCjjxqIfp1PqavH, ERpxhnx4yQO2gF4g0J9G8G, MDWW9wjzQsTkpJTsAXw1tG, OTCxoIqhEhA65VRuJvFoxB, PRVmCVU2hynJRxCDsjx8OE, a8xx20Fc5nKc8DbqSwNBuB, bPL0FcLvoxhO0amTUOV9QC, c1qRGYMEWodUPO7ZFq831QB, h7QHiA6jfRB0V5iS7nYrsR, l96dMLSJZGbzKOOaSawmDC, mgknRxAcgFrHqTt5CZvnSF, n65LdbEr6NMNaEFcjX8Fh6F, oFHbC0LQKaxvW8gPAQzBAB, pN9XTk8HB1jtfigsDxuKfE, r2jaHd7wMNX07DmqtoTGYfB, r4JngA0ZVhEElGRZci9fohF, sCFM4WicR6deeSAdSwumP, skXEjqLZnGZAr6RJ8QjjD, uUcj3UAzjmPW47yNyzbT8C, ucLx3e73qDSgpZETH1oJ9, uwZv0qzQLi0MDBWLWzKuAG, vLT6ef7BJliTDpt4k5jqF, w7JAMsElgYTLo8syEMZ8Lk, x9j7a5gok64zzNKnvdJNnE, yAfJq6fAufU3HOal8Q4DkG, yUuRVFmKCNYKHMIon8qCKG, yeHXFGHVMgEtZ4f1O7U2OB) begin U2JXBqjMcwW1AxVU5Q1ESG = ERpxhnx4yQO2gF4g0J9G8G; bm6UZNfjlfNI5cDV8oaTj = yAfJq6fAufU3HOal8Q4DkG; EzzigQlTGv8J7DBTRmqQ9C = yeHXFGHVMgEtZ4f1O7U2OB; srDEOQxwGboahrxQGs2vYE = w7JAMsElgYTLo8syEMZ8Lk; gZNZkxioohAMHXxms1BEOE = skXEjqLZnGZAr6RJ8QjjD; xhZyruBklMjVnVQHFCsnC = r2jaHd7wMNX07DmqtoTGYfB; MTuGLzs6sZnejyrpSaOMvF = MDWW9wjzQsTkpJTsAXw1tG; tArVqL2CTwuHoaoeSuZkaB = CDiyyho6hDs0nvcIRHvdfF; g4P4JTWbBBBn0JhReP8eXAH = EIQhCDitCjjxqIfp1PqavH; f1bIHzdG7kDHnL70sxnVWzB = PRVmCVU2hynJRxCDsjx8OE; s3m9T9rV2e4ZoMyZFS4lKeB = l96dMLSJZGbzKOOaSawmDC; p7ixx7ZWknoF1F7FbI5yjED = h7QHiA6jfRB0V5iS7nYrsR; KwC6wbRFLWpjZZERCcYIGB = pN9XTk8HB1jtfigsDxuKfE; MOh79n10Ewq3O8I6VYlcS = ucLx3e73qDSgpZETH1oJ9; Ym7Bnv0nBa8mPH5deUne6F = BAQ1YrOPn1tEt43kT1QPvE; e2MNnweVMUgzBGV1fQxq5dB = oFHbC0LQKaxvW8gPAQzBAB; A9eIucMmprrI3z0XPuKfq = yUuRVFmKCNYKHMIon8qCKG; CdyHxmDTkJd4Kce0MGL8uE = c1qRGYMEWodUPO7ZFq831QB; BlSFAnc8BhBCmuAIbP8voB = OTCxoIqhEhA65VRuJvFoxB; case ( oFHbC0LQKaxvW8gPAQzBAB) 3'b000 : begin s3m9T9rV2e4ZoMyZFS4lKeB = 16'sb0000000000000000; p7ixx7ZWknoF1F7FbI5yjED = 16'sb0000000000000000; KwC6wbRFLWpjZZERCcYIGB = 3'b000; Ym7Bnv0nBa8mPH5deUne6F = 3'b000; MOh79n10Ewq3O8I6VYlcS = 1'b0; BlSFAnc8BhBCmuAIbP8voB = 1'b0; e2MNnweVMUgzBGV1fQxq5dB = 3'b000; if ((c1qRGYMEWodUPO7ZFq831QB && (w7JAMsElgYTLo8syEMZ8Lk == 7'b1110111)) && PRVmCVU2hynJRxCDsjx8OE) begin s3m9T9rV2e4ZoMyZFS4lKeB = r4JngA0ZVhEElGRZci9fohF; p7ixx7ZWknoF1F7FbI5yjED = a8xx20Fc5nKc8DbqSwNBuB; KwC6wbRFLWpjZZERCcYIGB = 3'b000; if (vLT6ef7BJliTDpt4k5jqF) begin MOh79n10Ewq3O8I6VYlcS = 1'b1; e2MNnweVMUgzBGV1fQxq5dB = 3'b010; end else begin MOh79n10Ewq3O8I6VYlcS = 1'b0; e2MNnweVMUgzBGV1fQxq5dB = 3'b001; end end end 3'b001 : begin e2MNnweVMUgzBGV1fQxq5dB = 3'b001; BlSFAnc8BhBCmuAIbP8voB = 1'b0; if (vLT6ef7BJliTDpt4k5jqF) begin s3m9T9rV2e4ZoMyZFS4lKeB = r4JngA0ZVhEElGRZci9fohF; p7ixx7ZWknoF1F7FbI5yjED = a8xx20Fc5nKc8DbqSwNBuB; KwC6wbRFLWpjZZERCcYIGB = 3'b000; MOh79n10Ewq3O8I6VYlcS = 1'b1; e2MNnweVMUgzBGV1fQxq5dB = 3'b010; end end 3'b010 : begin s3m9T9rV2e4ZoMyZFS4lKeB = r4JngA0ZVhEElGRZci9fohF; p7ixx7ZWknoF1F7FbI5yjED = a8xx20Fc5nKc8DbqSwNBuB; BlSFAnc8BhBCmuAIbP8voB = 1'b0; if (pN9XTk8HB1jtfigsDxuKfE == 3'b111) begin MOh79n10Ewq3O8I6VYlcS = 1'b0; if (yUuRVFmKCNYKHMIon8qCKG) begin e2MNnweVMUgzBGV1fQxq5dB = 3'b100; BlSFAnc8BhBCmuAIbP8voB = 1'b1; Ym7Bnv0nBa8mPH5deUne6F = 3'b001; end else begin e2MNnweVMUgzBGV1fQxq5dB = 3'b011; end KwC6wbRFLWpjZZERCcYIGB = 3'b000; end else if (vLT6ef7BJliTDpt4k5jqF) begin e2MNnweVMUgzBGV1fQxq5dB = 3'b010; MOh79n10Ewq3O8I6VYlcS = 1'b1; KwC6wbRFLWpjZZERCcYIGB = pN9XTk8HB1jtfigsDxuKfE + 3'b001; end else begin e2MNnweVMUgzBGV1fQxq5dB = 3'b010; MOh79n10Ewq3O8I6VYlcS = 1'b0; end end 3'b011 : begin if (yUuRVFmKCNYKHMIon8qCKG) begin e2MNnweVMUgzBGV1fQxq5dB = 3'b100; BlSFAnc8BhBCmuAIbP8voB = 1'b1; Ym7Bnv0nBa8mPH5deUne6F = 3'b001; end end 3'b100 : begin if (BAQ1YrOPn1tEt43kT1QPvE == 3'b111) begin BlSFAnc8BhBCmuAIbP8voB = 1'b1; KwC6wbRFLWpjZZERCcYIGB = 3'b000; Ym7Bnv0nBa8mPH5deUne6F = 3'b000; if (c1qRGYMEWodUPO7ZFq831QB) begin s3m9T9rV2e4ZoMyZFS4lKeB = r4JngA0ZVhEElGRZci9fohF; p7ixx7ZWknoF1F7FbI5yjED = a8xx20Fc5nKc8DbqSwNBuB; if (vLT6ef7BJliTDpt4k5jqF) begin MOh79n10Ewq3O8I6VYlcS = 1'b1; e2MNnweVMUgzBGV1fQxq5dB = 3'b010; end else begin MOh79n10Ewq3O8I6VYlcS = 1'b0; e2MNnweVMUgzBGV1fQxq5dB = 3'b001; end end else begin e2MNnweVMUgzBGV1fQxq5dB = 3'b000; MOh79n10Ewq3O8I6VYlcS = 1'b0; s3m9T9rV2e4ZoMyZFS4lKeB = 16'sb0000000000000000; p7ixx7ZWknoF1F7FbI5yjED = 16'sb0000000000000000; end end else begin Ym7Bnv0nBa8mPH5deUne6F = BAQ1YrOPn1tEt43kT1QPvE + 3'b001; end end default : begin s3m9T9rV2e4ZoMyZFS4lKeB = 16'sb0000000000000000; p7ixx7ZWknoF1F7FbI5yjED = 16'sb0000000000000000; KwC6wbRFLWpjZZERCcYIGB = 3'b000; Ym7Bnv0nBa8mPH5deUne6F = 3'b000; MOh79n10Ewq3O8I6VYlcS = 1'b0; e2MNnweVMUgzBGV1fQxq5dB = 3'b000; end endcase case ( r2jaHd7wMNX07DmqtoTGYfB) 2'b00 : begin xhZyruBklMjVnVQHFCsnC = 2'b00; MTuGLzs6sZnejyrpSaOMvF = 7'b0000000; U2JXBqjMcwW1AxVU5Q1ESG = mgknRxAcgFrHqTt5CZvnSF; bm6UZNfjlfNI5cDV8oaTj = sCFM4WicR6deeSAdSwumP; EzzigQlTGv8J7DBTRmqQ9C = 1'b0; A9eIucMmprrI3z0XPuKfq = 1'b0; if (n65LdbEr6NMNaEFcjX8Fh6F) begin xhZyruBklMjVnVQHFCsnC = 2'b01; MTuGLzs6sZnejyrpSaOMvF = 7'b0000000; end end 2'b01 : begin xhZyruBklMjVnVQHFCsnC = 2'b01; A9eIucMmprrI3z0XPuKfq = 1'b0; if ((MDWW9wjzQsTkpJTsAXw1tG == 7'b1111111) && vLT6ef7BJliTDpt4k5jqF) begin xhZyruBklMjVnVQHFCsnC = 2'b10; end if (vLT6ef7BJliTDpt4k5jqF) begin MTuGLzs6sZnejyrpSaOMvF = MDWW9wjzQsTkpJTsAXw1tG + 7'b0000001; end U2JXBqjMcwW1AxVU5Q1ESG = x9j7a5gok64zzNKnvdJNnE; bm6UZNfjlfNI5cDV8oaTj = bPL0FcLvoxhO0amTUOV9QC; EzzigQlTGv8J7DBTRmqQ9C = vLT6ef7BJliTDpt4k5jqF; end 2'b10 : begin xhZyruBklMjVnVQHFCsnC = 2'b10; if ((MDWW9wjzQsTkpJTsAXw1tG == 7'b1110111) && BKNY6GzA6oGZumjzTATycD) begin xhZyruBklMjVnVQHFCsnC = 2'b01; A9eIucMmprrI3z0XPuKfq = 1'b1; end if (BKNY6GzA6oGZumjzTATycD) begin if (MDWW9wjzQsTkpJTsAXw1tG == 7'b1110111) begin MTuGLzs6sZnejyrpSaOMvF = 7'b0000000; end else begin MTuGLzs6sZnejyrpSaOMvF = MDWW9wjzQsTkpJTsAXw1tG + 7'b0000001; end end U2JXBqjMcwW1AxVU5Q1ESG = mgknRxAcgFrHqTt5CZvnSF; bm6UZNfjlfNI5cDV8oaTj = sCFM4WicR6deeSAdSwumP; EzzigQlTGv8J7DBTRmqQ9C = BKNY6GzA6oGZumjzTATycD; end default : begin xhZyruBklMjVnVQHFCsnC = 2'b00; MTuGLzs6sZnejyrpSaOMvF = 7'b0000000; U2JXBqjMcwW1AxVU5Q1ESG = mgknRxAcgFrHqTt5CZvnSF; bm6UZNfjlfNI5cDV8oaTj = sCFM4WicR6deeSAdSwumP; EzzigQlTGv8J7DBTRmqQ9C = BKNY6GzA6oGZumjzTATycD; end endcase case ( skXEjqLZnGZAr6RJ8QjjD) 3'b000 : begin gZNZkxioohAMHXxms1BEOE = 3'b000; CdyHxmDTkJd4Kce0MGL8uE = 1'b0; srDEOQxwGboahrxQGs2vYE = 7'b0000000; tArVqL2CTwuHoaoeSuZkaB = uUcj3UAzjmPW47yNyzbT8C; g4P4JTWbBBBn0JhReP8eXAH = uwZv0qzQLi0MDBWLWzKuAG; if (n65LdbEr6NMNaEFcjX8Fh6F) begin gZNZkxioohAMHXxms1BEOE = 3'b001; srDEOQxwGboahrxQGs2vYE = 7'b0000000; f1bIHzdG7kDHnL70sxnVWzB = 1'b1; end end 3'b001 : begin gZNZkxioohAMHXxms1BEOE = 3'b001; f1bIHzdG7kDHnL70sxnVWzB = 1'b0; CdyHxmDTkJd4Kce0MGL8uE = 1'b0; if (w7JAMsElgYTLo8syEMZ8Lk == 7'b1111111) begin if (vLT6ef7BJliTDpt4k5jqF) begin gZNZkxioohAMHXxms1BEOE = 3'b010; end else begin gZNZkxioohAMHXxms1BEOE = 3'b100; end srDEOQxwGboahrxQGs2vYE = 7'b0000000; f1bIHzdG7kDHnL70sxnVWzB = vLT6ef7BJliTDpt4k5jqF; tArVqL2CTwuHoaoeSuZkaB = r4JngA0ZVhEElGRZci9fohF; g4P4JTWbBBBn0JhReP8eXAH = a8xx20Fc5nKc8DbqSwNBuB; end else if (n65LdbEr6NMNaEFcjX8Fh6F) begin gZNZkxioohAMHXxms1BEOE = 3'b001; srDEOQxwGboahrxQGs2vYE = w7JAMsElgYTLo8syEMZ8Lk + 7'b0000001; f1bIHzdG7kDHnL70sxnVWzB = 1'b1; tArVqL2CTwuHoaoeSuZkaB = uUcj3UAzjmPW47yNyzbT8C; g4P4JTWbBBBn0JhReP8eXAH = uwZv0qzQLi0MDBWLWzKuAG; end end 3'b010 : begin gZNZkxioohAMHXxms1BEOE = 3'b010; f1bIHzdG7kDHnL70sxnVWzB = 1'b0; CdyHxmDTkJd4Kce0MGL8uE = 1'b0; if (w7JAMsElgYTLo8syEMZ8Lk == 7'b1110110) begin CdyHxmDTkJd4Kce0MGL8uE = 1'b1; end if (w7JAMsElgYTLo8syEMZ8Lk == 7'b1110111) begin srDEOQxwGboahrxQGs2vYE = w7JAMsElgYTLo8syEMZ8Lk + 7'b0000001; gZNZkxioohAMHXxms1BEOE = 3'b011; f1bIHzdG7kDHnL70sxnVWzB = 1'b0; tArVqL2CTwuHoaoeSuZkaB = uUcj3UAzjmPW47yNyzbT8C; g4P4JTWbBBBn0JhReP8eXAH = uwZv0qzQLi0MDBWLWzKuAG; end else if (vLT6ef7BJliTDpt4k5jqF) begin gZNZkxioohAMHXxms1BEOE = 3'b010; srDEOQxwGboahrxQGs2vYE = w7JAMsElgYTLo8syEMZ8Lk + 7'b0000001; f1bIHzdG7kDHnL70sxnVWzB = 1'b1; tArVqL2CTwuHoaoeSuZkaB = r4JngA0ZVhEElGRZci9fohF; g4P4JTWbBBBn0JhReP8eXAH = a8xx20Fc5nKc8DbqSwNBuB; end end 3'b011 : begin srDEOQxwGboahrxQGs2vYE = 7'b0000000; f1bIHzdG7kDHnL70sxnVWzB = n65LdbEr6NMNaEFcjX8Fh6F; tArVqL2CTwuHoaoeSuZkaB = uUcj3UAzjmPW47yNyzbT8C; g4P4JTWbBBBn0JhReP8eXAH = uwZv0qzQLi0MDBWLWzKuAG; CdyHxmDTkJd4Kce0MGL8uE = 1'b0; if (n65LdbEr6NMNaEFcjX8Fh6F) begin gZNZkxioohAMHXxms1BEOE = 3'b001; end else begin gZNZkxioohAMHXxms1BEOE = 3'b000; end end 3'b100 : begin gZNZkxioohAMHXxms1BEOE = 3'b100; f1bIHzdG7kDHnL70sxnVWzB = 1'b0; CdyHxmDTkJd4Kce0MGL8uE = 1'b0; if (vLT6ef7BJliTDpt4k5jqF) begin gZNZkxioohAMHXxms1BEOE = 3'b010; srDEOQxwGboahrxQGs2vYE = 7'b0000000; f1bIHzdG7kDHnL70sxnVWzB = 1'b1; tArVqL2CTwuHoaoeSuZkaB = r4JngA0ZVhEElGRZci9fohF; g4P4JTWbBBBn0JhReP8eXAH = a8xx20Fc5nKc8DbqSwNBuB; end end default : begin gZNZkxioohAMHXxms1BEOE = 3'b000; srDEOQxwGboahrxQGs2vYE = 7'b0000000; f1bIHzdG7kDHnL70sxnVWzB = n65LdbEr6NMNaEFcjX8Fh6F; tArVqL2CTwuHoaoeSuZkaB = uUcj3UAzjmPW47yNyzbT8C; g4P4JTWbBBBn0JhReP8eXAH = uwZv0qzQLi0MDBWLWzKuAG; end endcase r5kivPzvWgOSiA0gZBDsCMD = CDiyyho6hDs0nvcIRHvdfF; iOhy3XYM3su7ndksftfCZG = EIQhCDitCjjxqIfp1PqavH; TIIVgGzxbljXJKElx1RmZB = w7JAMsElgYTLo8syEMZ8Lk; d4GqKaFZXLUlts9HBCZPXG = PRVmCVU2hynJRxCDsjx8OE; lJc3nzBSuIub4Fgm41LhsH = l96dMLSJZGbzKOOaSawmDC; e4s7lktq7sxpTrarrx3LfPD = h7QHiA6jfRB0V5iS7nYrsR; mmaX8nGKzNYVdRyx6p1LtC = pN9XTk8HB1jtfigsDxuKfE; whMUFL1J2R7VsHTN9UxHOH = ucLx3e73qDSgpZETH1oJ9; pfAgd4CSuF40Tz4AXQRjjB = BAQ1YrOPn1tEt43kT1QPvE; tKu1I9axj5Jgdz0Uq0pTPF = OTCxoIqhEhA65VRuJvFoxB; rM5MTP4UKZC3il6lMwiHT = ERpxhnx4yQO2gF4g0J9G8G; gP6GlHEmSHKO19LfKcs3AH = yAfJq6fAufU3HOal8Q4DkG; wyxMTJhenZ0YDgDbHfiMlC = yeHXFGHVMgEtZ4f1O7U2OB; end PxGtD8RdpEuqNR1OqCny8D #(.AddrWidth(3), .DataWidth(16) ) t8AFKkvPqHL66Nrvwo08U3B (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .E7QNJoK4KvAThVFhUlvl2G(lJc3nzBSuIub4Fgm41LhsH), .l30d1QakAt61ivcMw8sJQE(mmaX8nGKzNYVdRyx6p1LtC), .UKo8akspo4h0jsZ6g712NB(whMUFL1J2R7VsHTN9UxHOH), .EYQG62ys4E6V8lISAdlW1C(pfAgd4CSuF40Tz4AXQRjjB), .HmVcl5yQin7hEovf3bwNG(PLGAQRVd1M1QgFrsMrWVBH) ); PxGtD8RdpEuqNR1OqCny8D #(.AddrWidth(3), .DataWidth(16) ) w0woCGNlGJrRwrjXj0Q0rC (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .E7QNJoK4KvAThVFhUlvl2G(e4s7lktq7sxpTrarrx3LfPD), .l30d1QakAt61ivcMw8sJQE(mmaX8nGKzNYVdRyx6p1LtC), .UKo8akspo4h0jsZ6g712NB(whMUFL1J2R7VsHTN9UxHOH), .EYQG62ys4E6V8lISAdlW1C(pfAgd4CSuF40Tz4AXQRjjB), .HmVcl5yQin7hEovf3bwNG(LifjwIUema6BHVuDJV77JF) ); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : f78KPhImpxKu3eA37uiPDC if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin cWUwraq7WjwtV5SP0dQobH <= 16'sb0000000000000000; v1iHIP96KWtHSOQsfIP0oDD <= 16'sb0000000000000000; r1RjufPwJY8CeBEsvwJ2flF <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin cWUwraq7WjwtV5SP0dQobH <= 16'sb0000000000000000; v1iHIP96KWtHSOQsfIP0oDD <= 16'sb0000000000000000; r1RjufPwJY8CeBEsvwJ2flF <= 1'b0; end else begin cWUwraq7WjwtV5SP0dQobH <= HVkI4mR4uVjbZBmf8GvOyF; v1iHIP96KWtHSOQsfIP0oDD <= VZmPcFtZLayUEhrt70JPkG; r1RjufPwJY8CeBEsvwJ2flF <= o59gL1lKXL2dKgQPA064uXG; end end end always @(LifjwIUema6BHVuDJV77JF, PLGAQRVd1M1QgFrsMrWVBH, cWUwraq7WjwtV5SP0dQobH, gP6GlHEmSHKO19LfKcs3AH, r1RjufPwJY8CeBEsvwJ2flF, rM5MTP4UKZC3il6lMwiHT, tKu1I9axj5Jgdz0Uq0pTPF, v1iHIP96KWtHSOQsfIP0oDD, wyxMTJhenZ0YDgDbHfiMlC) begin HVkI4mR4uVjbZBmf8GvOyF = cWUwraq7WjwtV5SP0dQobH; VZmPcFtZLayUEhrt70JPkG = v1iHIP96KWtHSOQsfIP0oDD; o59gL1lKXL2dKgQPA064uXG = r1RjufPwJY8CeBEsvwJ2flF; if (wyxMTJhenZ0YDgDbHfiMlC) begin HVkI4mR4uVjbZBmf8GvOyF = rM5MTP4UKZC3il6lMwiHT; VZmPcFtZLayUEhrt70JPkG = gP6GlHEmSHKO19LfKcs3AH; o59gL1lKXL2dKgQPA064uXG = 1'b1; end else if (tKu1I9axj5Jgdz0Uq0pTPF) begin HVkI4mR4uVjbZBmf8GvOyF = PLGAQRVd1M1QgFrsMrWVBH; VZmPcFtZLayUEhrt70JPkG = LifjwIUema6BHVuDJV77JF; o59gL1lKXL2dKgQPA064uXG = 1'b1; end else begin o59gL1lKXL2dKgQPA064uXG = 1'b0; end P3F2cuYaLRQxlfxwGBfSjF = cWUwraq7WjwtV5SP0dQobH; Rwrw0YN1HJLlhEzt1YbmaC = v1iHIP96KWtHSOQsfIP0oDD; vl2rwYFSlP59iBJIjf8F4D = r1RjufPwJY8CeBEsvwJ2flF; end assign N2ZdE4zLlq5uRV4rcE2wdE = r5kivPzvWgOSiA0gZBDsCMD; assign AECH0r3KnKo0RJFepDhYUD = TIIVgGzxbljXJKElx1RmZB; assign twcuYIJzeZMBjyHmZ1FZDD = d4GqKaFZXLUlts9HBCZPXG; assign f3NrgRvCkMfwf1E3PnKtczF = P3F2cuYaLRQxlfxwGBfSjF; assign f2XZKbXdctKWPTTQYeLkBWE = Rwrw0YN1HJLlhEzt1YbmaC; endmodule