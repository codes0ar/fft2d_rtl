`timescale 1 ns / 1 ns module PgyJIAY0PTIwvT911tPTDC (v04pHKxyc2sPW047bbyUgE, JAMOfrNHxGSYDF0urqkLN, l7IYN7joqiz566PVFOWVRgE, WJrLCpghLrgwyLgXr83JPE, gEaylbF1WXdCOYwXfvD4G, o4iXCc2GyRgQIsHmtR0i8nE, NdNevEoWljk83nSbsGDU1C, ymBdGOgDsRajoiY9d7TZdC, q8L6STCfvGEzwAAhXRTKviE, R6zf5iqRNVEGVBO8egq8kF, EnlAo7K66kKuzHIKWLmc1F, ew3EeLap6s8rXmNrsqaTWH, IPh1M0O3x0ioGlon72MROG, Mt05SNCQbo0cCPNa1yEFyF, Z7ZDy0EvwvoCh1zahAqvSF); input v04pHKxyc2sPW047bbyUgE; input JAMOfrNHxGSYDF0urqkLN; input signed [15:0] l7IYN7joqiz566PVFOWVRgE; input signed [15:0] WJrLCpghLrgwyLgXr83JPE; input signed [15:0] gEaylbF1WXdCOYwXfvD4G; input signed [15:0] o4iXCc2GyRgQIsHmtR0i8nE; input NdNevEoWljk83nSbsGDU1C; input signed [15:0] ymBdGOgDsRajoiY9d7TZdC; input signed [15:0] q8L6STCfvGEzwAAhXRTKviE; input R6zf5iqRNVEGVBO8egq8kF; output signed [15:0] EnlAo7K66kKuzHIKWLmc1F; output signed [15:0] ew3EeLap6s8rXmNrsqaTWH; output signed [15:0] IPh1M0O3x0ioGlon72MROG; output signed [15:0] Mt05SNCQbo0cCPNa1yEFyF; output Z7ZDy0EvwvoCh1zahAqvSF; reg signed [15:0] XOQBCWZyBA9fPc87mG5IsD; reg signed [15:0] jgpSuUOXE6beAUY2P4Iv4C; reg signed [15:0] s6mgKiePlUcVLouID5veYH; reg signed [15:0] Oze4Se7M5853Ky7frJBG9F; reg signed [15:0] MekY8xeaDEGsVWujfwtKYD; reg signed [15:0] umUHW18Nzczl7XvduT3KfG; reg signed [15:0] YhpEOQdmbC7NlFQDHpC9CG; reg signed [15:0] mHrFqLcAecA5gGbizXVkBB; reg signed [15:0] O2dufN5BaFwGqA9Oi3KkIC; reg signed [15:0] W3WuRCFnI5ngJZRPIZcluH; reg signed [15:0] PJ83Ne7TovKBk1QalAPkbF; reg signed [15:0] PQB4vyiY2hzUb277RaVY2G; reg signed [15:0] v1719E7mUU6xC7Ekf0pTEsD; reg signed [15:0] OAV4L8I57muqoGnQrH1vvB; reg signed [15:0] PYokxVN7N7QMAGDo8L7yrB; reg signed [15:0] t7SArk8uVG5hA9zEDrd2PB; reg signed [15:0] m5Y6o8AVvD1ar5547ejyQGD; reg signed [15:0] t5RODow4NCCeLJzE2dz9ImH; reg signed [15:0] Y4G0Jzpc0pu9WjWBN3cG3G; reg signed [15:0] yi5TBCH5TW5biX3U7QsRqE; reg signed [15:0] UV2a0iFkGBexVZbqWWEZtH; reg signed [15:0] srmdhX8C2dssNj53K6bvXB; reg signed [15:0] PI4X2832OFOysxpHuBiM9G; reg signed [15:0] wBO6oB2d6g6Z4IwDoFEshF; reg JRIoLUeCq9mXSVlgE57gFE; reg tSpBSFRas5hrgrmHKg0BzD; reg SNSO4dX03KiNOAsJChroeG; wire bV5IA5v0KhopEZ9ZLb20D; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : MczQYJ6MT1pYZD7C1UhQv if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin XOQBCWZyBA9fPc87mG5IsD <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin XOQBCWZyBA9fPc87mG5IsD <= 16'sb0000000000000000; end else begin XOQBCWZyBA9fPc87mG5IsD <= l7IYN7joqiz566PVFOWVRgE; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : xwyxj2YIc64Lxvl4r8S8mG if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin jgpSuUOXE6beAUY2P4Iv4C <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin jgpSuUOXE6beAUY2P4Iv4C <= 16'sb0000000000000000; end else begin jgpSuUOXE6beAUY2P4Iv4C <= XOQBCWZyBA9fPc87mG5IsD; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : L1HBH8O5DRbGBa9XvBX70C if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin s6mgKiePlUcVLouID5veYH <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin s6mgKiePlUcVLouID5veYH <= 16'sb0000000000000000; end else begin s6mgKiePlUcVLouID5veYH <= jgpSuUOXE6beAUY2P4Iv4C; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : s2CWr6rrksK4W7N0omU97HD if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin Oze4Se7M5853Ky7frJBG9F <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin Oze4Se7M5853Ky7frJBG9F <= 16'sb0000000000000000; end else begin Oze4Se7M5853Ky7frJBG9F <= s6mgKiePlUcVLouID5veYH; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : k1Zsi6BUVrSUjLbIYwh26G if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin MekY8xeaDEGsVWujfwtKYD <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin MekY8xeaDEGsVWujfwtKYD <= 16'sb0000000000000000; end else begin MekY8xeaDEGsVWujfwtKYD <= Oze4Se7M5853Ky7frJBG9F; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : TPi3Fu9uFLztbkFwa0H53D if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin umUHW18Nzczl7XvduT3KfG <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin umUHW18Nzczl7XvduT3KfG <= 16'sb0000000000000000; end else begin umUHW18Nzczl7XvduT3KfG <= MekY8xeaDEGsVWujfwtKYD; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : IBmSJmjQmOQZECy1AykU1D if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin YhpEOQdmbC7NlFQDHpC9CG <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin YhpEOQdmbC7NlFQDHpC9CG <= 16'sb0000000000000000; end else begin YhpEOQdmbC7NlFQDHpC9CG <= umUHW18Nzczl7XvduT3KfG; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : VNPcEW4KZxpAtEz0DCT8vD if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin mHrFqLcAecA5gGbizXVkBB <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin mHrFqLcAecA5gGbizXVkBB <= 16'sb0000000000000000; end else begin mHrFqLcAecA5gGbizXVkBB <= YhpEOQdmbC7NlFQDHpC9CG; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : t8uWAeIAh3IMbN9UNxoYBKD if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin O2dufN5BaFwGqA9Oi3KkIC <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin O2dufN5BaFwGqA9Oi3KkIC <= 16'sb0000000000000000; end else begin O2dufN5BaFwGqA9Oi3KkIC <= mHrFqLcAecA5gGbizXVkBB; end end end assign EnlAo7K66kKuzHIKWLmc1F = O2dufN5BaFwGqA9Oi3KkIC; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : QtzxgwI206U33aXvIkKdwD if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin W3WuRCFnI5ngJZRPIZcluH <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin W3WuRCFnI5ngJZRPIZcluH <= 16'sb0000000000000000; end else begin W3WuRCFnI5ngJZRPIZcluH <= WJrLCpghLrgwyLgXr83JPE; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : awX33YTQEl2OxkV2HHm04D if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin PJ83Ne7TovKBk1QalAPkbF <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin PJ83Ne7TovKBk1QalAPkbF <= 16'sb0000000000000000; end else begin PJ83Ne7TovKBk1QalAPkbF <= W3WuRCFnI5ngJZRPIZcluH; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : wroVmvZXsLz1H55Ur0PrpB if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin PQB4vyiY2hzUb277RaVY2G <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin PQB4vyiY2hzUb277RaVY2G <= 16'sb0000000000000000; end else begin PQB4vyiY2hzUb277RaVY2G <= PJ83Ne7TovKBk1QalAPkbF; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : z8NMcVNSFzdoHNpSsC5DBLF if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin v1719E7mUU6xC7Ekf0pTEsD <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin v1719E7mUU6xC7Ekf0pTEsD <= 16'sb0000000000000000; end else begin v1719E7mUU6xC7Ekf0pTEsD <= PQB4vyiY2hzUb277RaVY2G; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : j2gHN9roTaQcXLtCUWIL9F if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin OAV4L8I57muqoGnQrH1vvB <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin OAV4L8I57muqoGnQrH1vvB <= 16'sb0000000000000000; end else begin OAV4L8I57muqoGnQrH1vvB <= v1719E7mUU6xC7Ekf0pTEsD; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : eVDXDpbSTruDFXBM6ygPaB if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin PYokxVN7N7QMAGDo8L7yrB <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin PYokxVN7N7QMAGDo8L7yrB <= 16'sb0000000000000000; end else begin PYokxVN7N7QMAGDo8L7yrB <= OAV4L8I57muqoGnQrH1vvB; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : a2bprYW6bhaVvTUhwUfmVQF if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin t7SArk8uVG5hA9zEDrd2PB <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin t7SArk8uVG5hA9zEDrd2PB <= 16'sb0000000000000000; end else begin t7SArk8uVG5hA9zEDrd2PB <= PYokxVN7N7QMAGDo8L7yrB; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : RfFhiu7TcZArCuQWZZoVsB if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin m5Y6o8AVvD1ar5547ejyQGD <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin m5Y6o8AVvD1ar5547ejyQGD <= 16'sb0000000000000000; end else begin m5Y6o8AVvD1ar5547ejyQGD <= t7SArk8uVG5hA9zEDrd2PB; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : owLoaMKUokO7uUwJJovpJE if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin t5RODow4NCCeLJzE2dz9ImH <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin t5RODow4NCCeLJzE2dz9ImH <= 16'sb0000000000000000; end else begin t5RODow4NCCeLJzE2dz9ImH <= m5Y6o8AVvD1ar5547ejyQGD; end end end assign ew3EeLap6s8rXmNrsqaTWH = t5RODow4NCCeLJzE2dz9ImH; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : YKhHebQtfFPtGJB8AN9NfC if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin Y4G0Jzpc0pu9WjWBN3cG3G <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin Y4G0Jzpc0pu9WjWBN3cG3G <= 16'sb0000000000000000; end else begin Y4G0Jzpc0pu9WjWBN3cG3G <= gEaylbF1WXdCOYwXfvD4G; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : R02gF8dBxGuXtqNBiytOBD if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin yi5TBCH5TW5biX3U7QsRqE <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin yi5TBCH5TW5biX3U7QsRqE <= 16'sb0000000000000000; end else begin yi5TBCH5TW5biX3U7QsRqE <= Y4G0Jzpc0pu9WjWBN3cG3G; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : Fxt9eCqtG0jUXmLi6jZUvE if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin UV2a0iFkGBexVZbqWWEZtH <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin UV2a0iFkGBexVZbqWWEZtH <= 16'sb0000000000000000; end else begin UV2a0iFkGBexVZbqWWEZtH <= yi5TBCH5TW5biX3U7QsRqE; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : iRHyolisTvsKLxVejMexAB if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin srmdhX8C2dssNj53K6bvXB <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin srmdhX8C2dssNj53K6bvXB <= 16'sb0000000000000000; end else begin srmdhX8C2dssNj53K6bvXB <= o4iXCc2GyRgQIsHmtR0i8nE; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : e6AZe9KIcZJURxtpakQhtqG if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin PI4X2832OFOysxpHuBiM9G <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin PI4X2832OFOysxpHuBiM9G <= 16'sb0000000000000000; end else begin PI4X2832OFOysxpHuBiM9G <= srmdhX8C2dssNj53K6bvXB; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : y8LVueovJyghRSuIm8a5QH if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin wBO6oB2d6g6Z4IwDoFEshF <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin wBO6oB2d6g6Z4IwDoFEshF <= 16'sb0000000000000000; end else begin wBO6oB2d6g6Z4IwDoFEshF <= PI4X2832OFOysxpHuBiM9G; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : Yera4SjAVuKG7TjeL0xum if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin JRIoLUeCq9mXSVlgE57gFE <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin JRIoLUeCq9mXSVlgE57gFE <= 1'b0; end else begin JRIoLUeCq9mXSVlgE57gFE <= NdNevEoWljk83nSbsGDU1C; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : MplkH2AOPP4uw14V7wrk3B if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin tSpBSFRas5hrgrmHKg0BzD <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin tSpBSFRas5hrgrmHKg0BzD <= 1'b0; end else begin tSpBSFRas5hrgrmHKg0BzD <= JRIoLUeCq9mXSVlgE57gFE; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : QkTsAMX2ysQgjvkiAUs2oC if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin SNSO4dX03KiNOAsJChroeG <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin SNSO4dX03KiNOAsJChroeG <= 1'b0; end else begin SNSO4dX03KiNOAsJChroeG <= tSpBSFRas5hrgrmHKg0BzD; end end end GFWrW5VaXHBkOIv9SbevB JOQQNSibUv7LmaKv3pf63F (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .UV2a0iFkGBexVZbqWWEZtH(UV2a0iFkGBexVZbqWWEZtH), .wBO6oB2d6g6Z4IwDoFEshF(wBO6oB2d6g6Z4IwDoFEshF), .SNSO4dX03KiNOAsJChroeG(SNSO4dX03KiNOAsJChroeG), .ymBdGOgDsRajoiY9d7TZdC(ymBdGOgDsRajoiY9d7TZdC), .q8L6STCfvGEzwAAhXRTKviE(q8L6STCfvGEzwAAhXRTKviE), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .IPh1M0O3x0ioGlon72MROG(IPh1M0O3x0ioGlon72MROG), .Mt05SNCQbo0cCPNa1yEFyF(Mt05SNCQbo0cCPNa1yEFyF), .a3DgkQGhREeclbrZTuU8PBG(Z7ZDy0EvwvoCh1zahAqvSF) ); endmodule