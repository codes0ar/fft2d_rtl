`timescale 1 ns / 1 ns module uccCglqbDhsRCLPdxxn4OD (v04pHKxyc2sPW047bbyUgE, JAMOfrNHxGSYDF0urqkLN, lTYYhj3P59f6KeSXhObJAE, WawYOEnpsrkHlANz6YaiLG, l9QVSAqS6jsMaipvGnosLD, UwIsRF8C7ejj45D9sxKqgB, XVoYQfnVFtlWlmN3BG5OI, R6zf5iqRNVEGVBO8egq8kF, x3T5ivGGBQbBK8kZOoMj3, cMIOWiDVVCoNgM2IifcBEE, d7gCnTVLfOVVTEggcR6PDKC); input v04pHKxyc2sPW047bbyUgE; input JAMOfrNHxGSYDF0urqkLN; input signed [15:0] lTYYhj3P59f6KeSXhObJAE; input signed [15:0] WawYOEnpsrkHlANz6YaiLG; input l9QVSAqS6jsMaipvGnosLD; input signed [15:0] UwIsRF8C7ejj45D9sxKqgB; input signed [15:0] XVoYQfnVFtlWlmN3BG5OI; input R6zf5iqRNVEGVBO8egq8kF; output signed [15:0] x3T5ivGGBQbBK8kZOoMj3; output signed [15:0] cMIOWiDVVCoNgM2IifcBEE; output d7gCnTVLfOVVTEggcR6PDKC; reg signed [15:0] m8hJy2WxazSQVjwXAnlR7E; reg signed [15:0] TrIYqHGMr9KeALjla3ZjyF; reg signed [15:0] Qfqf2vuelr0iX7UmtewYhE; reg signed [15:0] n7GLhspJq27KHBdXHaZRPiE; reg signed [15:0] udARMRgYPzYB3bpLURr27B; reg signed [15:0] lqOJeKLhaKnwh3UOnSAeSG; reg signed [31:0] Pv40qULTbnH5xjOvV8bvvF; reg signed [31:0] xi6mK9xuygpCeLdYkgPJ2C; reg signed [31:0] CE2N9ZWS3erY7b120RyOSB; reg signed [31:0] x7XejrfM3CJ9nzMq4qWQClD; reg signed [15:0] aAj6KAvP6OSqCr33Vy4S1E; reg signed [15:0] pEfHnw2SW1hyYwjLZKqIv; reg signed [31:0] b8ky1cMhanM4yt6ecqpfeSD; reg signed [31:0] mhVUn1lDQRB9ezxqrc1oYE; reg signed [31:0] GRbpE81OwWRPPOX7uYPdCE; reg signed [31:0] ODjsec8sXmmf5oYetpkwF; reg l1dn5tWhZH93UlShOIFAV4C; reg zZkg29k58j3it2vW69T3rD; reg q7hX77ax2V3fGalwpJXdBH; reg nh1huyjuNrD92N6vFHOmDC; reg signed [32:0] y1QKCMUTAs3LMDFeQWvymFG; reg signed [32:0] h0vCcMropazUerM228ICNH; reg dd8BH6p2FEjlz6kiNafb5D; reg signed [31:0] V4BG2efg1IdmoaSGGxqsFB; reg signed [31:0] qX5r6geE6hwYyXsaJKR2VG; reg signed [31:0] pa8WlaH1GgDQDsT5FhgLPG; reg signed [31:0] MFPXFnqFXCXOmeBOqlKZ8C; wire signed [32:0] h5OyXxCHPUBY6X0KYzOKoE; wire signed [32:0] u3VKmh0jHfDtZBLwBdNHNR; wire signed [32:0] DX3ZtVdPStFPKnH25e2UHH; wire signed [32:0] v7rIbogJlhbqWkfHGbuGES; wire signed [32:0] r5BpjspgAgVeUPo7gCNUdC; wire signed [32:0] g7RI48YQk79hTwN3rQMThwD; wire signed [32:0] f2p28IFpladjvJgNAXEda5C; wire signed [32:0] pYqO0MCbB1ffrab9vhIynC; reg EJhGYSklU9oB2SMd4Kcpm; wire E8vXCbwD0Lvfu72APyVAvC; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : MczQYJ6MT1pYZD7C1UhQv if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin m8hJy2WxazSQVjwXAnlR7E <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin m8hJy2WxazSQVjwXAnlR7E <= 16'sb0000000000000000; end else begin m8hJy2WxazSQVjwXAnlR7E <= lTYYhj3P59f6KeSXhObJAE; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : xwyxj2YIc64Lxvl4r8S8mG if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin TrIYqHGMr9KeALjla3ZjyF <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin TrIYqHGMr9KeALjla3ZjyF <= 16'sb0000000000000000; end else begin TrIYqHGMr9KeALjla3ZjyF <= WawYOEnpsrkHlANz6YaiLG; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : L1HBH8O5DRbGBa9XvBX70C if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin Qfqf2vuelr0iX7UmtewYhE <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin Qfqf2vuelr0iX7UmtewYhE <= 16'sb0000000000000000; end else begin Qfqf2vuelr0iX7UmtewYhE <= UwIsRF8C7ejj45D9sxKqgB; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : s2CWr6rrksK4W7N0omU97HD if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin n7GLhspJq27KHBdXHaZRPiE <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin n7GLhspJq27KHBdXHaZRPiE <= 16'sb0000000000000000; end else begin n7GLhspJq27KHBdXHaZRPiE <= XVoYQfnVFtlWlmN3BG5OI; end end end always @(posedge v04pHKxyc2sPW047bbyUgE) begin : gbDxcjDe0CQuhiFjEnp8ED b8ky1cMhanM4yt6ecqpfeSD <= Pv40qULTbnH5xjOvV8bvvF; GRbpE81OwWRPPOX7uYPdCE <= xi6mK9xuygpCeLdYkgPJ2C; mhVUn1lDQRB9ezxqrc1oYE <= CE2N9ZWS3erY7b120RyOSB; ODjsec8sXmmf5oYetpkwF <= x7XejrfM3CJ9nzMq4qWQClD; Pv40qULTbnH5xjOvV8bvvF <= udARMRgYPzYB3bpLURr27B * aAj6KAvP6OSqCr33Vy4S1E; xi6mK9xuygpCeLdYkgPJ2C <= lqOJeKLhaKnwh3UOnSAeSG * pEfHnw2SW1hyYwjLZKqIv; CE2N9ZWS3erY7b120RyOSB <= udARMRgYPzYB3bpLURr27B * pEfHnw2SW1hyYwjLZKqIv; x7XejrfM3CJ9nzMq4qWQClD <= lqOJeKLhaKnwh3UOnSAeSG * aAj6KAvP6OSqCr33Vy4S1E; aAj6KAvP6OSqCr33Vy4S1E <= Qfqf2vuelr0iX7UmtewYhE; pEfHnw2SW1hyYwjLZKqIv <= n7GLhspJq27KHBdXHaZRPiE; udARMRgYPzYB3bpLURr27B <= m8hJy2WxazSQVjwXAnlR7E; lqOJeKLhaKnwh3UOnSAeSG <= TrIYqHGMr9KeALjla3ZjyF; end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : k1Zsi6BUVrSUjLbIYwh26G if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin l1dn5tWhZH93UlShOIFAV4C <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin l1dn5tWhZH93UlShOIFAV4C <= 1'b0; end else begin l1dn5tWhZH93UlShOIFAV4C <= l9QVSAqS6jsMaipvGnosLD; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : TPi3Fu9uFLztbkFwa0H53D if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin zZkg29k58j3it2vW69T3rD <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin zZkg29k58j3it2vW69T3rD <= 1'b0; end else begin zZkg29k58j3it2vW69T3rD <= l1dn5tWhZH93UlShOIFAV4C; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : IBmSJmjQmOQZECy1AykU1D if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin q7hX77ax2V3fGalwpJXdBH <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin q7hX77ax2V3fGalwpJXdBH <= 1'b0; end else begin q7hX77ax2V3fGalwpJXdBH <= zZkg29k58j3it2vW69T3rD; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : VNPcEW4KZxpAtEz0DCT8vD if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin nh1huyjuNrD92N6vFHOmDC <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin nh1huyjuNrD92N6vFHOmDC <= 1'b0; end else begin nh1huyjuNrD92N6vFHOmDC <= q7hX77ax2V3fGalwpJXdBH; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : P4xI0OA7WlHTOpYREhqff if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin y1QKCMUTAs3LMDFeQWvymFG <= 33'sh000000000; h0vCcMropazUerM228ICNH <= 33'sh000000000; V4BG2efg1IdmoaSGGxqsFB <= 32'sb00000000000000000000000000000000; qX5r6geE6hwYyXsaJKR2VG <= 32'sb00000000000000000000000000000000; pa8WlaH1GgDQDsT5FhgLPG <= 32'sb00000000000000000000000000000000; MFPXFnqFXCXOmeBOqlKZ8C <= 32'sb00000000000000000000000000000000; dd8BH6p2FEjlz6kiNafb5D <= 1'b0; EJhGYSklU9oB2SMd4Kcpm <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin y1QKCMUTAs3LMDFeQWvymFG <= 33'sh000000000; h0vCcMropazUerM228ICNH <= 33'sh000000000; V4BG2efg1IdmoaSGGxqsFB <= 32'sb00000000000000000000000000000000; qX5r6geE6hwYyXsaJKR2VG <= 32'sb00000000000000000000000000000000; pa8WlaH1GgDQDsT5FhgLPG <= 32'sb00000000000000000000000000000000; MFPXFnqFXCXOmeBOqlKZ8C <= 32'sb00000000000000000000000000000000; dd8BH6p2FEjlz6kiNafb5D <= 1'b0; EJhGYSklU9oB2SMd4Kcpm <= 1'b0; end else begin y1QKCMUTAs3LMDFeQWvymFG <= h5OyXxCHPUBY6X0KYzOKoE; h0vCcMropazUerM228ICNH <= u3VKmh0jHfDtZBLwBdNHNR; V4BG2efg1IdmoaSGGxqsFB <= b8ky1cMhanM4yt6ecqpfeSD; qX5r6geE6hwYyXsaJKR2VG <= mhVUn1lDQRB9ezxqrc1oYE; pa8WlaH1GgDQDsT5FhgLPG <= GRbpE81OwWRPPOX7uYPdCE; MFPXFnqFXCXOmeBOqlKZ8C <= ODjsec8sXmmf5oYetpkwF; EJhGYSklU9oB2SMd4Kcpm <= dd8BH6p2FEjlz6kiNafb5D; dd8BH6p2FEjlz6kiNafb5D <= nh1huyjuNrD92N6vFHOmDC; end end end assign DX3ZtVdPStFPKnH25e2UHH = {V4BG2efg1IdmoaSGGxqsFB[31], V4BG2efg1IdmoaSGGxqsFB}; assign v7rIbogJlhbqWkfHGbuGES = {pa8WlaH1GgDQDsT5FhgLPG[31], pa8WlaH1GgDQDsT5FhgLPG}; assign h5OyXxCHPUBY6X0KYzOKoE = DX3ZtVdPStFPKnH25e2UHH - v7rIbogJlhbqWkfHGbuGES; assign r5BpjspgAgVeUPo7gCNUdC = {qX5r6geE6hwYyXsaJKR2VG[31], qX5r6geE6hwYyXsaJKR2VG}; assign g7RI48YQk79hTwN3rQMThwD = {MFPXFnqFXCXOmeBOqlKZ8C[31], MFPXFnqFXCXOmeBOqlKZ8C}; assign u3VKmh0jHfDtZBLwBdNHNR = r5BpjspgAgVeUPo7gCNUdC + g7RI48YQk79hTwN3rQMThwD; assign f2p28IFpladjvJgNAXEda5C = y1QKCMUTAs3LMDFeQWvymFG; assign pYqO0MCbB1ffrab9vhIynC = h0vCcMropazUerM228ICNH; assign x3T5ivGGBQbBK8kZOoMj3 = f2p28IFpladjvJgNAXEda5C[29:14] + $signed({1'b0, f2p28IFpladjvJgNAXEda5C[13]}); assign cMIOWiDVVCoNgM2IifcBEE = pYqO0MCbB1ffrab9vhIynC[29:14] + $signed({1'b0, pYqO0MCbB1ffrab9vhIynC[13]}); assign d7gCnTVLfOVVTEggcR6PDKC = EJhGYSklU9oB2SMd4Kcpm; endmodule