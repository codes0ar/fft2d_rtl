`timescale 1 ns / 1 ns module q2kRA8XOHHRNcp89kCO6bC (v04pHKxyc2sPW047bbyUgE, JAMOfrNHxGSYDF0urqkLN, Pq4nKEqqr18aLXK1kX1dfH, R6zf5iqRNVEGVBO8egq8kF, mvb8xVo6CcFPFyQu3ctDE, gC05dypmmuscVux3EfDHCD); input v04pHKxyc2sPW047bbyUgE; input JAMOfrNHxGSYDF0urqkLN; input Pq4nKEqqr18aLXK1kX1dfH; input R6zf5iqRNVEGVBO8egq8kF; output signed [15:0] mvb8xVo6CcFPFyQu3ctDE; output signed [15:0] gC05dypmmuscVux3EfDHCD; reg [4:0] TE2s9kaW4jbT2yuidpcUIF; reg [1:0] j9GInQQXHbUGPAy0R0X4BQD; reg [2:0] URO3uEJ9VVi4n2rv5pG4XF; reg [6:0] mevVutOyAH9CPJEBvvvxsF; reg [3:0] Mndh5cWFT2MK7irxEkUgvB; reg DSwbuqNl6si2qBBlHlS4m; reg ADYssd29ifP9Cnqtxk4KFH; reg zUwvjmWVganUujWHX9Ik8G; reg [4:0] vyYw1SbJbcSwGlwsC50cRF; reg [1:0] tHBJR87iWmyApKoUBwoC; reg [2:0] ZXzEhgRyMkDiwOKQ1ZyHtH; reg [6:0] vndcJtBZasetzBa7iOZamH; reg [3:0] W3LV4fQGt3vLDwUnzRRUwH; reg t96JNxh4AbzBXPo2zT29dlG; reg ARo3kgZ8gBa9Exsckya1UB; reg IvvfGB2My0fbqvU6mi859D; reg [3:0] DOFNWCpbdQSLsWtzwny1qG; reg EWvO8Kf2QN2SS53GJJcWwF; reg [2:0] j9HNozHmNa6lYL8HVho1pB; reg B9qRWWVXUMKaf08lKjOj5G; wire signed [15:0] zVla2Vy8BUCugJ5Gig2ZK [0:15]; wire signed [15:0] F8NQxbAEqqIEtFo6mesHd; reg signed [15:0] CIRDDBHrGgCpm7HNrbXUCF; wire signed [15:0] ysWUViVY5R4DChvjvp5gDD [0:15]; wire signed [15:0] jsn1oqDToTuWwgUlIvqN3; reg signed [15:0] M9MMs7oRisnNmiBXjmtOsD; reg [2:0] YjlT6Mg9KMpPzxF47HzV7D; reg UrNpVdQvuAmKReKH4NECKD; reg signed [15:0] ONIgquJLgLedZU10qrtlZG; reg signed [15:0] Tcw9zGJiOCDLQO3MwcKjnC; reg [2:0] CbpoQEK97vFu56nv3223yC; reg [6:0] xouA8rA79zSw8rxilmdIcF; reg [4:0] GW0FC9j2OjlJb11BmqyTwH; reg signed [15:0] uCEkpKGKs7tQvr2GeEGSGC; reg signed [15:0] hhzTcPgpleSJBYLOoujKGG; reg signed [8:0] cVX5EXK4yxLZ1cYzNgyXx; reg signed [8:0] g4zMZYWhK020aMvVlufXSO; reg signed [15:0] SVYTAuHmM7AdeQD3dklB3D; reg signed [15:0] z9uPanlNUawhpWBfZzoV6C; reg signed [15:0] iKPA1JOFbNoLsuo87UbsvD; reg signed [15:0] K3fvtqFABfYnMEzDvYIrq; reg signed [8:0] jbCFxKpbanHjkeuxNFuv1D; reg signed [8:0] xs6NJDxbN0KSgBeqxxDWYF; reg signed [15:0] KwiyVhhhZdTrDQCbiLV8zE; reg signed [15:0] sGNGvuvL8Q7LZvZSVKC57B; reg signed [16:0] WJY0hyRMua5sU8DuMmLu4; reg signed [16:0] b6ofl8SS59auHuq7NOO0WOG; reg signed [16:0] f2RPd8CpcTyQnKsmtWEywG; reg signed [16:0] w4sUCJ8sn9dqukS5aRJDigE; reg signed [16:0] L3USkDc1T9xpZF6CkNG03D; reg signed [16:0] s195ulFHSeSTCYTLhumIdD; wire VgCXfMa1NOcWXjwcxjhVAG; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : A7mAa8MkEw1SBVJbtTHnZE if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin URO3uEJ9VVi4n2rv5pG4XF <= 3'b000; mevVutOyAH9CPJEBvvvxsF <= 7'b0000000; Mndh5cWFT2MK7irxEkUgvB <= 4'b0000; DSwbuqNl6si2qBBlHlS4m <= 1'b0; ADYssd29ifP9Cnqtxk4KFH <= 1'b0; zUwvjmWVganUujWHX9Ik8G <= 1'b0; TE2s9kaW4jbT2yuidpcUIF <= 5'b00000; j9GInQQXHbUGPAy0R0X4BQD <= 2'b11; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin URO3uEJ9VVi4n2rv5pG4XF <= 3'b000; mevVutOyAH9CPJEBvvvxsF <= 7'b0000000; Mndh5cWFT2MK7irxEkUgvB <= 4'b0000; DSwbuqNl6si2qBBlHlS4m <= 1'b0; ADYssd29ifP9Cnqtxk4KFH <= 1'b0; zUwvjmWVganUujWHX9Ik8G <= 1'b0; TE2s9kaW4jbT2yuidpcUIF <= 5'b00000; j9GInQQXHbUGPAy0R0X4BQD <= 2'b11; end else begin TE2s9kaW4jbT2yuidpcUIF <= vyYw1SbJbcSwGlwsC50cRF; j9GInQQXHbUGPAy0R0X4BQD <= tHBJR87iWmyApKoUBwoC; URO3uEJ9VVi4n2rv5pG4XF <= ZXzEhgRyMkDiwOKQ1ZyHtH; mevVutOyAH9CPJEBvvvxsF <= vndcJtBZasetzBa7iOZamH; Mndh5cWFT2MK7irxEkUgvB <= W3LV4fQGt3vLDwUnzRRUwH; DSwbuqNl6si2qBBlHlS4m <= t96JNxh4AbzBXPo2zT29dlG; ADYssd29ifP9Cnqtxk4KFH <= ARo3kgZ8gBa9Exsckya1UB; zUwvjmWVganUujWHX9Ik8G <= IvvfGB2My0fbqvU6mi859D; end end end always @(ADYssd29ifP9Cnqtxk4KFH, DSwbuqNl6si2qBBlHlS4m, Mndh5cWFT2MK7irxEkUgvB, Pq4nKEqqr18aLXK1kX1dfH, TE2s9kaW4jbT2yuidpcUIF, URO3uEJ9VVi4n2rv5pG4XF, j9GInQQXHbUGPAy0R0X4BQD, mevVutOyAH9CPJEBvvvxsF, zUwvjmWVganUujWHX9Ik8G) begin hhzTcPgpleSJBYLOoujKGG = 16'sb0000000000000000; cVX5EXK4yxLZ1cYzNgyXx = 9'sb000000000; g4zMZYWhK020aMvVlufXSO = 9'sb000000000; z9uPanlNUawhpWBfZzoV6C = 16'sb0000000000000000; K3fvtqFABfYnMEzDvYIrq = 16'sb0000000000000000; xouA8rA79zSw8rxilmdIcF = 7'b0000000; uCEkpKGKs7tQvr2GeEGSGC = 16'sb0000000000000000; SVYTAuHmM7AdeQD3dklB3D = 16'sb0000000000000000; iKPA1JOFbNoLsuo87UbsvD = 16'sb0000000000000000; jbCFxKpbanHjkeuxNFuv1D = 9'sb000000000; xs6NJDxbN0KSgBeqxxDWYF = 9'sb000000000; vyYw1SbJbcSwGlwsC50cRF = TE2s9kaW4jbT2yuidpcUIF; tHBJR87iWmyApKoUBwoC = j9GInQQXHbUGPAy0R0X4BQD; vndcJtBZasetzBa7iOZamH = mevVutOyAH9CPJEBvvvxsF; W3LV4fQGt3vLDwUnzRRUwH = Mndh5cWFT2MK7irxEkUgvB; t96JNxh4AbzBXPo2zT29dlG = DSwbuqNl6si2qBBlHlS4m; IvvfGB2My0fbqvU6mi859D = ADYssd29ifP9Cnqtxk4KFH; ARo3kgZ8gBa9Exsckya1UB = Pq4nKEqqr18aLXK1kX1dfH; case ( mevVutOyAH9CPJEBvvvxsF) 7'b0010000 : begin CbpoQEK97vFu56nv3223yC = 3'b000; t96JNxh4AbzBXPo2zT29dlG = 1'b1; end 7'b0100000 : begin CbpoQEK97vFu56nv3223yC = 3'b001; t96JNxh4AbzBXPo2zT29dlG = 1'b0; end 7'b0110000 : begin CbpoQEK97vFu56nv3223yC = 3'b010; t96JNxh4AbzBXPo2zT29dlG = 1'b1; end 7'b1000000 : begin CbpoQEK97vFu56nv3223yC = 3'b011; t96JNxh4AbzBXPo2zT29dlG = 1'b0; end 7'b1010000 : begin CbpoQEK97vFu56nv3223yC = 3'b100; t96JNxh4AbzBXPo2zT29dlG = 1'b1; end default : begin CbpoQEK97vFu56nv3223yC = mevVutOyAH9CPJEBvvvxsF[6:4]; t96JNxh4AbzBXPo2zT29dlG = 1'b0; end endcase ZXzEhgRyMkDiwOKQ1ZyHtH = CbpoQEK97vFu56nv3223yC; case ( CbpoQEK97vFu56nv3223yC) 3'b000 : begin W3LV4fQGt3vLDwUnzRRUwH = mevVutOyAH9CPJEBvvvxsF[3:0]; end 3'b001 : begin jbCFxKpbanHjkeuxNFuv1D = {2'b0, mevVutOyAH9CPJEBvvvxsF}; cVX5EXK4yxLZ1cYzNgyXx = 9'sb000100000 - jbCFxKpbanHjkeuxNFuv1D; W3LV4fQGt3vLDwUnzRRUwH = cVX5EXK4yxLZ1cYzNgyXx[3:0]; end 3'b010 : begin xs6NJDxbN0KSgBeqxxDWYF = {2'b0, mevVutOyAH9CPJEBvvvxsF}; g4zMZYWhK020aMvVlufXSO = xs6NJDxbN0KSgBeqxxDWYF - 9'sb000100000; W3LV4fQGt3vLDwUnzRRUwH = g4zMZYWhK020aMvVlufXSO[3:0]; end 3'b011 : begin SVYTAuHmM7AdeQD3dklB3D = {5'b0, {mevVutOyAH9CPJEBvvvxsF, 4'b0000}}; z9uPanlNUawhpWBfZzoV6C = 16'sb0000010000000000 - SVYTAuHmM7AdeQD3dklB3D; W3LV4fQGt3vLDwUnzRRUwH = z9uPanlNUawhpWBfZzoV6C[7:4]; end 3'b100 : begin iKPA1JOFbNoLsuo87UbsvD = {5'b0, {mevVutOyAH9CPJEBvvvxsF, 4'b0000}}; K3fvtqFABfYnMEzDvYIrq = iKPA1JOFbNoLsuo87UbsvD - 16'sb0000010000000000; W3LV4fQGt3vLDwUnzRRUwH = K3fvtqFABfYnMEzDvYIrq[7:4]; end default : begin uCEkpKGKs7tQvr2GeEGSGC = {5'b0, {mevVutOyAH9CPJEBvvvxsF, 4'b0000}}; hhzTcPgpleSJBYLOoujKGG = 16'sb0000011000000000 - uCEkpKGKs7tQvr2GeEGSGC; W3LV4fQGt3vLDwUnzRRUwH = hhzTcPgpleSJBYLOoujKGG[7:4]; end endcase GW0FC9j2OjlJb11BmqyTwH = {TE2s9kaW4jbT2yuidpcUIF[0], TE2s9kaW4jbT2yuidpcUIF[1], TE2s9kaW4jbT2yuidpcUIF[2], TE2s9kaW4jbT2yuidpcUIF[3], TE2s9kaW4jbT2yuidpcUIF[4]}; if (j9GInQQXHbUGPAy0R0X4BQD == 2'b00) begin vndcJtBZasetzBa7iOZamH = 7'b0000000; end else if (j9GInQQXHbUGPAy0R0X4BQD == 2'b01) begin vndcJtBZasetzBa7iOZamH = {2'b0, GW0FC9j2OjlJb11BmqyTwH}; end else if (j9GInQQXHbUGPAy0R0X4BQD == 2'b10) begin vndcJtBZasetzBa7iOZamH = {2'b0, GW0FC9j2OjlJb11BmqyTwH} <<< 8'd1; end else begin xouA8rA79zSw8rxilmdIcF = {2'b0, GW0FC9j2OjlJb11BmqyTwH}; vndcJtBZasetzBa7iOZamH = (xouA8rA79zSw8rxilmdIcF <<< 8'd1) + xouA8rA79zSw8rxilmdIcF; end if (Pq4nKEqqr18aLXK1kX1dfH) begin vyYw1SbJbcSwGlwsC50cRF = TE2s9kaW4jbT2yuidpcUIF + 5'b00001; end DOFNWCpbdQSLsWtzwny1qG = Mndh5cWFT2MK7irxEkUgvB; EWvO8Kf2QN2SS53GJJcWwF = zUwvjmWVganUujWHX9Ik8G; j9HNozHmNa6lYL8HVho1pB = URO3uEJ9VVi4n2rv5pG4XF; B9qRWWVXUMKaf08lKjOj5G = DSwbuqNl6si2qBBlHlS4m; end assign zVla2Vy8BUCugJ5Gig2ZK[0] = 16'sb0100000000000000; assign zVla2Vy8BUCugJ5Gig2ZK[1] = 16'sb0011111111101100; assign zVla2Vy8BUCugJ5Gig2ZK[2] = 16'sb0011111110110001; assign zVla2Vy8BUCugJ5Gig2ZK[3] = 16'sb0011111101001111; assign zVla2Vy8BUCugJ5Gig2ZK[4] = 16'sb0011111011000101; assign zVla2Vy8BUCugJ5Gig2ZK[5] = 16'sb0011111000010101; assign zVla2Vy8BUCugJ5Gig2ZK[6] = 16'sb0011110100111111; assign zVla2Vy8BUCugJ5Gig2ZK[7] = 16'sb0011110001000010; assign zVla2Vy8BUCugJ5Gig2ZK[8] = 16'sb0011101100100001; assign zVla2Vy8BUCugJ5Gig2ZK[9] = 16'sb0011100111011011; assign zVla2Vy8BUCugJ5Gig2ZK[10] = 16'sb0011100001110001; assign zVla2Vy8BUCugJ5Gig2ZK[11] = 16'sb0011011011100101; assign zVla2Vy8BUCugJ5Gig2ZK[12] = 16'sb0011010100110111; assign zVla2Vy8BUCugJ5Gig2ZK[13] = 16'sb0011001101101000; assign zVla2Vy8BUCugJ5Gig2ZK[14] = 16'sb0011000101111001; assign zVla2Vy8BUCugJ5Gig2ZK[15] = 16'sb0010111101101100; assign F8NQxbAEqqIEtFo6mesHd = zVla2Vy8BUCugJ5Gig2ZK[DOFNWCpbdQSLsWtzwny1qG]; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : j0boDGRQkCezKyDxbtKinG if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin CIRDDBHrGgCpm7HNrbXUCF <= 16'sb0000000000000000; end else begin CIRDDBHrGgCpm7HNrbXUCF <= F8NQxbAEqqIEtFo6mesHd; end end assign ysWUViVY5R4DChvjvp5gDD[0] = 16'sb0000000000000000; assign ysWUViVY5R4DChvjvp5gDD[1] = 16'sb1111110011011100; assign ysWUViVY5R4DChvjvp5gDD[2] = 16'sb1111100110111010; assign ysWUViVY5R4DChvjvp5gDD[3] = 16'sb1111011010011100; assign ysWUViVY5R4DChvjvp5gDD[4] = 16'sb1111001110000100; assign ysWUViVY5R4DChvjvp5gDD[5] = 16'sb1111000001110011; assign ysWUViVY5R4DChvjvp5gDD[6] = 16'sb1110110101101100; assign ysWUViVY5R4DChvjvp5gDD[7] = 16'sb1110101001110000; assign ysWUViVY5R4DChvjvp5gDD[8] = 16'sb1110011110000010; assign ysWUViVY5R4DChvjvp5gDD[9] = 16'sb1110010010100011; assign ysWUViVY5R4DChvjvp5gDD[10] = 16'sb1110000111010101; assign ysWUViVY5R4DChvjvp5gDD[11] = 16'sb1101111100011001; assign ysWUViVY5R4DChvjvp5gDD[12] = 16'sb1101110001110010; assign ysWUViVY5R4DChvjvp5gDD[13] = 16'sb1101100111100000; assign ysWUViVY5R4DChvjvp5gDD[14] = 16'sb1101011101100110; assign ysWUViVY5R4DChvjvp5gDD[15] = 16'sb1101010100000101; assign jsn1oqDToTuWwgUlIvqN3 = ysWUViVY5R4DChvjvp5gDD[DOFNWCpbdQSLsWtzwny1qG]; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : VAVA4twBRLX2WfwOrbR5l if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin M9MMs7oRisnNmiBXjmtOsD <= 16'sb0000000000000000; end else begin M9MMs7oRisnNmiBXjmtOsD <= jsn1oqDToTuWwgUlIvqN3; end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : MczQYJ6MT1pYZD7C1UhQv if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin YjlT6Mg9KMpPzxF47HzV7D <= 3'b000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin YjlT6Mg9KMpPzxF47HzV7D <= 3'b000; end else begin YjlT6Mg9KMpPzxF47HzV7D <= j9HNozHmNa6lYL8HVho1pB; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : xwyxj2YIc64Lxvl4r8S8mG if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin UrNpVdQvuAmKReKH4NECKD <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin UrNpVdQvuAmKReKH4NECKD <= 1'b0; end else begin UrNpVdQvuAmKReKH4NECKD <= B9qRWWVXUMKaf08lKjOj5G; end end end always @(CIRDDBHrGgCpm7HNrbXUCF, M9MMs7oRisnNmiBXjmtOsD, UrNpVdQvuAmKReKH4NECKD, YjlT6Mg9KMpPzxF47HzV7D) begin WJY0hyRMua5sU8DuMmLu4 = 17'sb00000000000000000; b6ofl8SS59auHuq7NOO0WOG = 17'sb00000000000000000; f2RPd8CpcTyQnKsmtWEywG = 17'sb00000000000000000; w4sUCJ8sn9dqukS5aRJDigE = 17'sb00000000000000000; L3USkDc1T9xpZF6CkNG03D = 17'sb00000000000000000; s195ulFHSeSTCYTLhumIdD = 17'sb00000000000000000; KwiyVhhhZdTrDQCbiLV8zE = CIRDDBHrGgCpm7HNrbXUCF; sGNGvuvL8Q7LZvZSVKC57B = M9MMs7oRisnNmiBXjmtOsD; if (UrNpVdQvuAmKReKH4NECKD) begin case ( YjlT6Mg9KMpPzxF47HzV7D) 3'b000 : begin KwiyVhhhZdTrDQCbiLV8zE = 16'sb0010110101000001; sGNGvuvL8Q7LZvZSVKC57B = 16'sb1101001010111111; end 3'b010 : begin KwiyVhhhZdTrDQCbiLV8zE = 16'sb1101001010111111; sGNGvuvL8Q7LZvZSVKC57B = 16'sb1101001010111111; end 3'b100 : begin KwiyVhhhZdTrDQCbiLV8zE = 16'sb1101001010111111; sGNGvuvL8Q7LZvZSVKC57B = 16'sb0010110101000001; end default : begin KwiyVhhhZdTrDQCbiLV8zE = 16'sb0010110101000001; sGNGvuvL8Q7LZvZSVKC57B = 16'sb1101001010111111; end endcase end else begin case ( YjlT6Mg9KMpPzxF47HzV7D) 3'b000 : begin end 3'b001 : begin WJY0hyRMua5sU8DuMmLu4 = - ({M9MMs7oRisnNmiBXjmtOsD[15], M9MMs7oRisnNmiBXjmtOsD}); KwiyVhhhZdTrDQCbiLV8zE = WJY0hyRMua5sU8DuMmLu4[15:0]; w4sUCJ8sn9dqukS5aRJDigE = - ({CIRDDBHrGgCpm7HNrbXUCF[15], CIRDDBHrGgCpm7HNrbXUCF}); sGNGvuvL8Q7LZvZSVKC57B = w4sUCJ8sn9dqukS5aRJDigE[15:0]; end 3'b010 : begin KwiyVhhhZdTrDQCbiLV8zE = M9MMs7oRisnNmiBXjmtOsD; L3USkDc1T9xpZF6CkNG03D = - ({CIRDDBHrGgCpm7HNrbXUCF[15], CIRDDBHrGgCpm7HNrbXUCF}); sGNGvuvL8Q7LZvZSVKC57B = L3USkDc1T9xpZF6CkNG03D[15:0]; end 3'b011 : begin b6ofl8SS59auHuq7NOO0WOG = - ({CIRDDBHrGgCpm7HNrbXUCF[15], CIRDDBHrGgCpm7HNrbXUCF}); KwiyVhhhZdTrDQCbiLV8zE = b6ofl8SS59auHuq7NOO0WOG[15:0]; sGNGvuvL8Q7LZvZSVKC57B = M9MMs7oRisnNmiBXjmtOsD; end 3'b100 : begin f2RPd8CpcTyQnKsmtWEywG = - ({CIRDDBHrGgCpm7HNrbXUCF[15], CIRDDBHrGgCpm7HNrbXUCF}); KwiyVhhhZdTrDQCbiLV8zE = f2RPd8CpcTyQnKsmtWEywG[15:0]; s195ulFHSeSTCYTLhumIdD = - ({M9MMs7oRisnNmiBXjmtOsD[15], M9MMs7oRisnNmiBXjmtOsD}); sGNGvuvL8Q7LZvZSVKC57B = s195ulFHSeSTCYTLhumIdD[15:0]; end default : begin KwiyVhhhZdTrDQCbiLV8zE = M9MMs7oRisnNmiBXjmtOsD; sGNGvuvL8Q7LZvZSVKC57B = CIRDDBHrGgCpm7HNrbXUCF; end endcase end ONIgquJLgLedZU10qrtlZG = KwiyVhhhZdTrDQCbiLV8zE; Tcw9zGJiOCDLQO3MwcKjnC = sGNGvuvL8Q7LZvZSVKC57B; end assign mvb8xVo6CcFPFyQu3ctDE = ONIgquJLgLedZU10qrtlZG; assign gC05dypmmuscVux3EfDHCD = Tcw9zGJiOCDLQO3MwcKjnC; endmodule