`timescale 1 ns / 1 ns module yp36yVdBki2iBRVFYzbmt (v04pHKxyc2sPW047bbyUgE, JAMOfrNHxGSYDF0urqkLN, EIYK1nT0oJLxbcxjmodwrC, l45qCeMpWMHOXjwYLaHORRE, j8SzfGJHmeoXnV9bhAUk40F, dMKGmQc7XAB1i3kk2Yk0hH, ydI2XfENb2Kl0A3qJMSMBB, nXMdpgmOgBwUAR30aQsd0B, kenMGol9N3qu644VwSIQzD, ovgS7leqdS5z2NH8xqTyeH, eWSF2FqZGP4L33XPl3WfqF, KgtpP4p0xLhni3stSN9j2F, bcPgddVda1xlzyptajDlFG, kUUVLVsgipRk0xKvCGrGvE); input v04pHKxyc2sPW047bbyUgE; input JAMOfrNHxGSYDF0urqkLN; input signed [15:0] EIYK1nT0oJLxbcxjmodwrC; input signed [15:0] l45qCeMpWMHOXjwYLaHORRE; input signed [15:0] j8SzfGJHmeoXnV9bhAUk40F; input signed [15:0] dMKGmQc7XAB1i3kk2Yk0hH; input signed [15:0] ydI2XfENb2Kl0A3qJMSMBB; input signed [15:0] nXMdpgmOgBwUAR30aQsd0B; input signed [15:0] kenMGol9N3qu644VwSIQzD; input signed [15:0] ovgS7leqdS5z2NH8xqTyeH; output [15:0] eWSF2FqZGP4L33XPl3WfqF; output [15:0] KgtpP4p0xLhni3stSN9j2F; output [15:0] bcPgddVda1xlzyptajDlFG; output [15:0] kUUVLVsgipRk0xKvCGrGvE; wire signed [15:0] sxjBgfCPJWPEwO3RfuCJLF [0:3]; wire signed [31:0] ZQPBCaH3CsAL98Ma7SQotB [0:3]; wire signed [15:0] ENys1xr2aw310RHqQ3zdZH [0:3]; wire signed [31:0] n1itWMDc2h5j1fFOw38UqmH [0:3]; wire [31:0] l7diY0oAQ4WZLEHmxtcnKl; wire [31:0] LoEbG9xSpCVNUBMqr4b6m; wire [32:0] lFIFc1FMCEhdqlYwYW5oSD; wire [31:0] ILjRXb7j5xUya5k8e6PTwD; wire [31:0] bZpzmZ2GtI3INKevWSVlzC; wire [32:0] DB14wLF62mIfBaTI6vec6B; wire [31:0] H20cUpLhsfVfJ92LJAQOWD; wire [31:0] jwMQr349SzDWq73ix7hnt; wire [32:0] DdWFbmNZw3i61r2Flc3lJG; wire [31:0] xLdGXDAP9TpO5keaXtpUCE; wire [31:0] NUZ0cOiLhQfqUrn215R0iF; wire [32:0] x2qOSwxaMdgo7eci0FxvvcF; wire [31:0] vuZ2nTtiQpIZLJSUSetjMF [0:3]; wire [15:0] waa48Uw91SZFWZY9mU7nvC; wire [15:0] ZO8mjpSGYWl4VDPzeaquoG; wire [15:0] kw2ymNvc9MOkxm4Ou30fqB; wire [15:0] BolOGJJauVSqkQjNqvMtlD; wire c54WqZL42iYdnhuPevgzcvC; assign sxjBgfCPJWPEwO3RfuCJLF[0] = EIYK1nT0oJLxbcxjmodwrC; assign sxjBgfCPJWPEwO3RfuCJLF[1] = l45qCeMpWMHOXjwYLaHORRE; assign sxjBgfCPJWPEwO3RfuCJLF[2] = j8SzfGJHmeoXnV9bhAUk40F; assign sxjBgfCPJWPEwO3RfuCJLF[3] = dMKGmQc7XAB1i3kk2Yk0hH; assign ZQPBCaH3CsAL98Ma7SQotB[0] = sxjBgfCPJWPEwO3RfuCJLF[0] * sxjBgfCPJWPEwO3RfuCJLF[0]; assign ZQPBCaH3CsAL98Ma7SQotB[1] = sxjBgfCPJWPEwO3RfuCJLF[1] * sxjBgfCPJWPEwO3RfuCJLF[1]; assign ZQPBCaH3CsAL98Ma7SQotB[2] = sxjBgfCPJWPEwO3RfuCJLF[2] * sxjBgfCPJWPEwO3RfuCJLF[2]; assign ZQPBCaH3CsAL98Ma7SQotB[3] = sxjBgfCPJWPEwO3RfuCJLF[3] * sxjBgfCPJWPEwO3RfuCJLF[3]; assign ENys1xr2aw310RHqQ3zdZH[0] = ydI2XfENb2Kl0A3qJMSMBB; assign ENys1xr2aw310RHqQ3zdZH[1] = nXMdpgmOgBwUAR30aQsd0B; assign ENys1xr2aw310RHqQ3zdZH[2] = kenMGol9N3qu644VwSIQzD; assign ENys1xr2aw310RHqQ3zdZH[3] = ovgS7leqdS5z2NH8xqTyeH; assign n1itWMDc2h5j1fFOw38UqmH[0] = ENys1xr2aw310RHqQ3zdZH[0] * ENys1xr2aw310RHqQ3zdZH[0]; assign n1itWMDc2h5j1fFOw38UqmH[1] = ENys1xr2aw310RHqQ3zdZH[1] * ENys1xr2aw310RHqQ3zdZH[1]; assign n1itWMDc2h5j1fFOw38UqmH[2] = ENys1xr2aw310RHqQ3zdZH[2] * ENys1xr2aw310RHqQ3zdZH[2]; assign n1itWMDc2h5j1fFOw38UqmH[3] = ENys1xr2aw310RHqQ3zdZH[3] * ENys1xr2aw310RHqQ3zdZH[3]; assign l7diY0oAQ4WZLEHmxtcnKl = (ZQPBCaH3CsAL98Ma7SQotB[0][31] == 1'b1 ? 32'b00000000000000000000000000000000 : ZQPBCaH3CsAL98Ma7SQotB[0]); assign LoEbG9xSpCVNUBMqr4b6m = (n1itWMDc2h5j1fFOw38UqmH[0][31] == 1'b1 ? 32'b00000000000000000000000000000000 : n1itWMDc2h5j1fFOw38UqmH[0]); assign lFIFc1FMCEhdqlYwYW5oSD = ({1'b0, l7diY0oAQ4WZLEHmxtcnKl}) + ({1'b0, LoEbG9xSpCVNUBMqr4b6m}); assign vuZ2nTtiQpIZLJSUSetjMF[0] = (lFIFc1FMCEhdqlYwYW5oSD[32] != 1'b0 ? 32'b11111111111111111111111111111111 : lFIFc1FMCEhdqlYwYW5oSD[31:0]); assign ILjRXb7j5xUya5k8e6PTwD = (ZQPBCaH3CsAL98Ma7SQotB[1][31] == 1'b1 ? 32'b00000000000000000000000000000000 : ZQPBCaH3CsAL98Ma7SQotB[1]); assign bZpzmZ2GtI3INKevWSVlzC = (n1itWMDc2h5j1fFOw38UqmH[1][31] == 1'b1 ? 32'b00000000000000000000000000000000 : n1itWMDc2h5j1fFOw38UqmH[1]); assign DB14wLF62mIfBaTI6vec6B = ({1'b0, ILjRXb7j5xUya5k8e6PTwD}) + ({1'b0, bZpzmZ2GtI3INKevWSVlzC}); assign vuZ2nTtiQpIZLJSUSetjMF[1] = (DB14wLF62mIfBaTI6vec6B[32] != 1'b0 ? 32'b11111111111111111111111111111111 : DB14wLF62mIfBaTI6vec6B[31:0]); assign H20cUpLhsfVfJ92LJAQOWD = (ZQPBCaH3CsAL98Ma7SQotB[2][31] == 1'b1 ? 32'b00000000000000000000000000000000 : ZQPBCaH3CsAL98Ma7SQotB[2]); assign jwMQr349SzDWq73ix7hnt = (n1itWMDc2h5j1fFOw38UqmH[2][31] == 1'b1 ? 32'b00000000000000000000000000000000 : n1itWMDc2h5j1fFOw38UqmH[2]); assign DdWFbmNZw3i61r2Flc3lJG = ({1'b0, H20cUpLhsfVfJ92LJAQOWD}) + ({1'b0, jwMQr349SzDWq73ix7hnt}); assign vuZ2nTtiQpIZLJSUSetjMF[2] = (DdWFbmNZw3i61r2Flc3lJG[32] != 1'b0 ? 32'b11111111111111111111111111111111 : DdWFbmNZw3i61r2Flc3lJG[31:0]); assign xLdGXDAP9TpO5keaXtpUCE = (ZQPBCaH3CsAL98Ma7SQotB[3][31] == 1'b1 ? 32'b00000000000000000000000000000000 : ZQPBCaH3CsAL98Ma7SQotB[3]); assign NUZ0cOiLhQfqUrn215R0iF = (n1itWMDc2h5j1fFOw38UqmH[3][31] == 1'b1 ? 32'b00000000000000000000000000000000 : n1itWMDc2h5j1fFOw38UqmH[3]); assign x2qOSwxaMdgo7eci0FxvvcF = ({1'b0, xLdGXDAP9TpO5keaXtpUCE}) + ({1'b0, NUZ0cOiLhQfqUrn215R0iF}); assign vuZ2nTtiQpIZLJSUSetjMF[3] = (x2qOSwxaMdgo7eci0FxvvcF[32] != 1'b0 ? 32'b11111111111111111111111111111111 : x2qOSwxaMdgo7eci0FxvvcF[31:0]); IWIdafyrOBWRPUGK17dNTF l4y2MZWq6Aps8DsHv33WzBC (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .h4h0SDZC9CQgXKPbimISL3(vuZ2nTtiQpIZLJSUSetjMF[0]), .b0pPxQrhAhYENzTiTGGny5G(vuZ2nTtiQpIZLJSUSetjMF[1]), .jQKNLtXo0Dqi6Vn3Jy2niG(vuZ2nTtiQpIZLJSUSetjMF[2]), .rosLsgtHKD6hJ64eM2pegF(vuZ2nTtiQpIZLJSUSetjMF[3]), .j71O4t3Nm1w5MRqcbOUNtHF(waa48Uw91SZFWZY9mU7nvC), .DVmjaezJpTmh9E1RX58vDE(ZO8mjpSGYWl4VDPzeaquoG), .c50jzfprXP85SKSfjge64NC(kw2ymNvc9MOkxm4Ou30fqB), .s7ASYYS329kRVgP7KY37Y(BolOGJJauVSqkQjNqvMtlD) ); assign eWSF2FqZGP4L33XPl3WfqF = waa48Uw91SZFWZY9mU7nvC; assign KgtpP4p0xLhni3stSN9j2F = ZO8mjpSGYWl4VDPzeaquoG; assign bcPgddVda1xlzyptajDlFG = kw2ymNvc9MOkxm4Ou30fqB; assign kUUVLVsgipRk0xKvCGrGvE = BolOGJJauVSqkQjNqvMtlD; endmodule