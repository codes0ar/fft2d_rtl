`timescale 1 ns / 1 ns module rUdEDJxz9hCFSCEPZfs0dH (v04pHKxyc2sPW047bbyUgE, JAMOfrNHxGSYDF0urqkLN, QWAACQosHJOUrDgm1wJeoG, hKoHLVfoAgFN4AYEXJutV, R6zf5iqRNVEGVBO8egq8kF, WgU2KCxd1j6m3EUCPiuf1F, y9Hu20tqKGzmg7O1xqeuAZH, F9FfK0xrG2zVVJqYJzgfxD, xGMN0H1JXsbMHEVz1iuteB); input v04pHKxyc2sPW047bbyUgE; input JAMOfrNHxGSYDF0urqkLN; input QWAACQosHJOUrDgm1wJeoG; input hKoHLVfoAgFN4AYEXJutV; input R6zf5iqRNVEGVBO8egq8kF; output WgU2KCxd1j6m3EUCPiuf1F; output y9Hu20tqKGzmg7O1xqeuAZH; output F9FfK0xrG2zVVJqYJzgfxD; output xGMN0H1JXsbMHEVz1iuteB; reg [1:0] X7FJ0jgk6hqdMN8BingGvE; reg [1:0] WXS42gmgDxS46057b3AGD; reg GP01IUV0xObQQCSdqL463C; reg [1:0] mb13NdjIe7rpJDLNih8AaE; reg [1:0] xSW8arCNXsyV5zIEXuGUQB; reg [1:0] ck9Ya76HU61qWvvl3qwfRG; reg dQhJtS5aSGZCPWaJqkkHi; reg [1:0] BNI9VucWF1TWsCAM4sBCHE; reg leyi2m0N7tcSGqQt5ZuKiH; reg o7vmW4wfrdqol0SHVeNyjHF; reg fEO4OYnhf0Uvi4JmepMxfB; reg vYfyltvUNNiXC2DaoA0A3F; wire i9zNkMcI7ViljEiLkC2zRjH; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : h6oTzWU1a3otHwaiji95ID if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin GP01IUV0xObQQCSdqL463C <= 1'b0; X7FJ0jgk6hqdMN8BingGvE <= 2'b00; WXS42gmgDxS46057b3AGD <= 2'b00; mb13NdjIe7rpJDLNih8AaE <= 2'b00; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin GP01IUV0xObQQCSdqL463C <= 1'b0; X7FJ0jgk6hqdMN8BingGvE <= 2'b00; WXS42gmgDxS46057b3AGD <= 2'b00; mb13NdjIe7rpJDLNih8AaE <= 2'b00; end else begin X7FJ0jgk6hqdMN8BingGvE <= xSW8arCNXsyV5zIEXuGUQB; WXS42gmgDxS46057b3AGD <= ck9Ya76HU61qWvvl3qwfRG; GP01IUV0xObQQCSdqL463C <= dQhJtS5aSGZCPWaJqkkHi; mb13NdjIe7rpJDLNih8AaE <= BNI9VucWF1TWsCAM4sBCHE; end end end always @(GP01IUV0xObQQCSdqL463C, QWAACQosHJOUrDgm1wJeoG, WXS42gmgDxS46057b3AGD, X7FJ0jgk6hqdMN8BingGvE, hKoHLVfoAgFN4AYEXJutV, mb13NdjIe7rpJDLNih8AaE) begin xSW8arCNXsyV5zIEXuGUQB = X7FJ0jgk6hqdMN8BingGvE; ck9Ya76HU61qWvvl3qwfRG = WXS42gmgDxS46057b3AGD; dQhJtS5aSGZCPWaJqkkHi = GP01IUV0xObQQCSdqL463C; BNI9VucWF1TWsCAM4sBCHE = mb13NdjIe7rpJDLNih8AaE; case ( mb13NdjIe7rpJDLNih8AaE) 2'b00 : begin BNI9VucWF1TWsCAM4sBCHE = 2'b00; vYfyltvUNNiXC2DaoA0A3F = 1'b0; if (WXS42gmgDxS46057b3AGD == 2'b01) begin BNI9VucWF1TWsCAM4sBCHE = 2'b01; end end 2'b01 : begin vYfyltvUNNiXC2DaoA0A3F = 1'b0; if (WXS42gmgDxS46057b3AGD == 2'b00) begin BNI9VucWF1TWsCAM4sBCHE = 2'b10; end end 2'b10 : begin vYfyltvUNNiXC2DaoA0A3F = 1'b0; BNI9VucWF1TWsCAM4sBCHE = 2'b11; end 2'b11 : begin vYfyltvUNNiXC2DaoA0A3F = 1'b1; BNI9VucWF1TWsCAM4sBCHE = 2'b00; end default : begin BNI9VucWF1TWsCAM4sBCHE = 2'b00; vYfyltvUNNiXC2DaoA0A3F = 1'b0; end endcase case ( WXS42gmgDxS46057b3AGD) 2'b00 : begin ck9Ya76HU61qWvvl3qwfRG = 2'b00; dQhJtS5aSGZCPWaJqkkHi = 1'b0; o7vmW4wfrdqol0SHVeNyjHF = 1'b0; if ((X7FJ0jgk6hqdMN8BingGvE == 2'b11) && QWAACQosHJOUrDgm1wJeoG) begin ck9Ya76HU61qWvvl3qwfRG = 2'b01; o7vmW4wfrdqol0SHVeNyjHF = hKoHLVfoAgFN4AYEXJutV; end end 2'b01 : begin o7vmW4wfrdqol0SHVeNyjHF = hKoHLVfoAgFN4AYEXJutV; if (hKoHLVfoAgFN4AYEXJutV) begin ck9Ya76HU61qWvvl3qwfRG = 2'b00; end end default : begin ck9Ya76HU61qWvvl3qwfRG = 2'b00; dQhJtS5aSGZCPWaJqkkHi = 1'b0; o7vmW4wfrdqol0SHVeNyjHF = 1'b0; end endcase case ( X7FJ0jgk6hqdMN8BingGvE) 2'b00 : begin xSW8arCNXsyV5zIEXuGUQB = 2'b00; fEO4OYnhf0Uvi4JmepMxfB = 1'b0; if (QWAACQosHJOUrDgm1wJeoG) begin xSW8arCNXsyV5zIEXuGUQB = 2'b11; end end 2'b11 : begin xSW8arCNXsyV5zIEXuGUQB = 2'b11; fEO4OYnhf0Uvi4JmepMxfB = 1'b0; if (QWAACQosHJOUrDgm1wJeoG) begin xSW8arCNXsyV5zIEXuGUQB = 2'b10; fEO4OYnhf0Uvi4JmepMxfB = 1'b1; end end 2'b10 : begin fEO4OYnhf0Uvi4JmepMxfB = 1'b0; xSW8arCNXsyV5zIEXuGUQB = 2'b10; if (QWAACQosHJOUrDgm1wJeoG) begin xSW8arCNXsyV5zIEXuGUQB = 2'b11; end end default : begin xSW8arCNXsyV5zIEXuGUQB = 2'b00; fEO4OYnhf0Uvi4JmepMxfB = 1'b0; end endcase leyi2m0N7tcSGqQt5ZuKiH = GP01IUV0xObQQCSdqL463C; end assign WgU2KCxd1j6m3EUCPiuf1F = leyi2m0N7tcSGqQt5ZuKiH; assign y9Hu20tqKGzmg7O1xqeuAZH = o7vmW4wfrdqol0SHVeNyjHF; assign F9FfK0xrG2zVVJqYJzgfxD = fEO4OYnhf0Uvi4JmepMxfB; assign xGMN0H1JXsbMHEVz1iuteB = vYfyltvUNNiXC2DaoA0A3F; endmodule