`timescale 1 ns / 1 ns module CQ8VhzX2aZDdqpzcRKBClF (v04pHKxyc2sPW047bbyUgE, JAMOfrNHxGSYDF0urqkLN, m0Pt9awzMYrRUb1BRHcMLqG, o3XsAkfAYoavjVukPhwjwlC, R6zf5iqRNVEGVBO8egq8kF, g1oJwDFAtNAcPvLahTlMEB, wf5f4XnltnQYt1bEDWEp0F, Q7D2KKVRLkwEPktPhyCkSD); input v04pHKxyc2sPW047bbyUgE; input JAMOfrNHxGSYDF0urqkLN; input m0Pt9awzMYrRUb1BRHcMLqG; input o3XsAkfAYoavjVukPhwjwlC; input R6zf5iqRNVEGVBO8egq8kF; output g1oJwDFAtNAcPvLahTlMEB; output wf5f4XnltnQYt1bEDWEp0F; output Q7D2KKVRLkwEPktPhyCkSD; reg JomiEQo6ylRrlhLJPFsQTG; reg [1:0] X7FJ0jgk6hqdMN8BingGvE; reg [1:0] WXS42gmgDxS46057b3AGD; reg GP01IUV0xObQQCSdqL463C; reg pDYTWTp6fyrEdA1XnDiP6E; reg [1:0] mb13NdjIe7rpJDLNih8AaE; reg Xf88wK4mkniJ6qfkmOXy2C; reg i2IIQfdSjOGJ0HAlaZdYe; reg [1:0] xSW8arCNXsyV5zIEXuGUQB; reg [1:0] ck9Ya76HU61qWvvl3qwfRG; reg dQhJtS5aSGZCPWaJqkkHi; reg t69iUVjqBKXZw2tNuE5YceG; reg [1:0] BNI9VucWF1TWsCAM4sBCHE; reg EIfu64RX7LMQGnynQeCGuD; reg euwYuFBjOyzJ1StMM7x9lB; reg n40UqkH7P32znVloyhHzXD; reg qhMTHhfDKHqjrVnmTgdY6; reg pBYDq5TsLLci7qFUEEbLfB; wire Qypqp0u3orfGM435LYgoJF; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : h6oTzWU1a3otHwaiji95ID if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin JomiEQo6ylRrlhLJPFsQTG <= 1'b0; GP01IUV0xObQQCSdqL463C <= 1'b0; X7FJ0jgk6hqdMN8BingGvE <= 2'b00; WXS42gmgDxS46057b3AGD <= 2'b00; mb13NdjIe7rpJDLNih8AaE <= 2'b00; pDYTWTp6fyrEdA1XnDiP6E <= 1'b0; Xf88wK4mkniJ6qfkmOXy2C <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin JomiEQo6ylRrlhLJPFsQTG <= 1'b0; GP01IUV0xObQQCSdqL463C <= 1'b0; X7FJ0jgk6hqdMN8BingGvE <= 2'b00; WXS42gmgDxS46057b3AGD <= 2'b00; mb13NdjIe7rpJDLNih8AaE <= 2'b00; pDYTWTp6fyrEdA1XnDiP6E <= 1'b0; Xf88wK4mkniJ6qfkmOXy2C <= 1'b0; end else begin JomiEQo6ylRrlhLJPFsQTG <= i2IIQfdSjOGJ0HAlaZdYe; X7FJ0jgk6hqdMN8BingGvE <= xSW8arCNXsyV5zIEXuGUQB; WXS42gmgDxS46057b3AGD <= ck9Ya76HU61qWvvl3qwfRG; GP01IUV0xObQQCSdqL463C <= dQhJtS5aSGZCPWaJqkkHi; pDYTWTp6fyrEdA1XnDiP6E <= t69iUVjqBKXZw2tNuE5YceG; mb13NdjIe7rpJDLNih8AaE <= BNI9VucWF1TWsCAM4sBCHE; Xf88wK4mkniJ6qfkmOXy2C <= EIfu64RX7LMQGnynQeCGuD; end end end always @(GP01IUV0xObQQCSdqL463C, JomiEQo6ylRrlhLJPFsQTG, WXS42gmgDxS46057b3AGD, X7FJ0jgk6hqdMN8BingGvE, Xf88wK4mkniJ6qfkmOXy2C, m0Pt9awzMYrRUb1BRHcMLqG, mb13NdjIe7rpJDLNih8AaE, o3XsAkfAYoavjVukPhwjwlC, pDYTWTp6fyrEdA1XnDiP6E) begin i2IIQfdSjOGJ0HAlaZdYe = JomiEQo6ylRrlhLJPFsQTG; xSW8arCNXsyV5zIEXuGUQB = X7FJ0jgk6hqdMN8BingGvE; ck9Ya76HU61qWvvl3qwfRG = WXS42gmgDxS46057b3AGD; dQhJtS5aSGZCPWaJqkkHi = GP01IUV0xObQQCSdqL463C; t69iUVjqBKXZw2tNuE5YceG = pDYTWTp6fyrEdA1XnDiP6E; BNI9VucWF1TWsCAM4sBCHE = mb13NdjIe7rpJDLNih8AaE; EIfu64RX7LMQGnynQeCGuD = Xf88wK4mkniJ6qfkmOXy2C; case ( mb13NdjIe7rpJDLNih8AaE) 2'b00 : begin BNI9VucWF1TWsCAM4sBCHE = 2'b00; EIfu64RX7LMQGnynQeCGuD = 1'b0; if (WXS42gmgDxS46057b3AGD == 2'b01) begin BNI9VucWF1TWsCAM4sBCHE = 2'b01; end end 2'b01 : begin EIfu64RX7LMQGnynQeCGuD = 1'b0; if (WXS42gmgDxS46057b3AGD == 2'b10) begin BNI9VucWF1TWsCAM4sBCHE = 2'b10; end end 2'b10 : begin EIfu64RX7LMQGnynQeCGuD = 1'b0; if (WXS42gmgDxS46057b3AGD == 2'b01) begin BNI9VucWF1TWsCAM4sBCHE = 2'b11; EIfu64RX7LMQGnynQeCGuD = 1'b1; end end 2'b11 : begin if (WXS42gmgDxS46057b3AGD == 2'b01) begin BNI9VucWF1TWsCAM4sBCHE = 2'b11; EIfu64RX7LMQGnynQeCGuD = 1'b1; end else begin EIfu64RX7LMQGnynQeCGuD = 1'b0; BNI9VucWF1TWsCAM4sBCHE = 2'b00; end end default : begin BNI9VucWF1TWsCAM4sBCHE = 2'b00; EIfu64RX7LMQGnynQeCGuD = 1'b0; end endcase case ( WXS42gmgDxS46057b3AGD) 2'b00 : begin ck9Ya76HU61qWvvl3qwfRG = 2'b00; dQhJtS5aSGZCPWaJqkkHi = 1'b0; n40UqkH7P32znVloyhHzXD = 1'b0; if (pDYTWTp6fyrEdA1XnDiP6E) begin ck9Ya76HU61qWvvl3qwfRG = 2'b01; n40UqkH7P32znVloyhHzXD = o3XsAkfAYoavjVukPhwjwlC; if (o3XsAkfAYoavjVukPhwjwlC) begin dQhJtS5aSGZCPWaJqkkHi = 1'b1; end end end 2'b01 : begin ck9Ya76HU61qWvvl3qwfRG = 2'b01; n40UqkH7P32znVloyhHzXD = o3XsAkfAYoavjVukPhwjwlC; if (o3XsAkfAYoavjVukPhwjwlC) begin if (GP01IUV0xObQQCSdqL463C == 1'b1) begin ck9Ya76HU61qWvvl3qwfRG = 2'b10; dQhJtS5aSGZCPWaJqkkHi = 1'b0; end else begin dQhJtS5aSGZCPWaJqkkHi = 1'b1; end end end 2'b10 : begin n40UqkH7P32znVloyhHzXD = 1'b0; if (GP01IUV0xObQQCSdqL463C == 1'b1) begin dQhJtS5aSGZCPWaJqkkHi = 1'b0; if (pDYTWTp6fyrEdA1XnDiP6E) begin ck9Ya76HU61qWvvl3qwfRG = 2'b01; end else begin ck9Ya76HU61qWvvl3qwfRG = 2'b00; end end else begin dQhJtS5aSGZCPWaJqkkHi = 1'b1; end end default : begin ck9Ya76HU61qWvvl3qwfRG = 2'b00; dQhJtS5aSGZCPWaJqkkHi = 1'b0; n40UqkH7P32znVloyhHzXD = 1'b0; end endcase case ( X7FJ0jgk6hqdMN8BingGvE) 2'b00 : begin xSW8arCNXsyV5zIEXuGUQB = 2'b00; i2IIQfdSjOGJ0HAlaZdYe = 1'b0; t69iUVjqBKXZw2tNuE5YceG = 1'b0; if (m0Pt9awzMYrRUb1BRHcMLqG) begin xSW8arCNXsyV5zIEXuGUQB = 2'b01; i2IIQfdSjOGJ0HAlaZdYe = 1'b1; end end 2'b01 : begin xSW8arCNXsyV5zIEXuGUQB = 2'b01; t69iUVjqBKXZw2tNuE5YceG = 1'b0; if (m0Pt9awzMYrRUb1BRHcMLqG) begin xSW8arCNXsyV5zIEXuGUQB = 2'b10; t69iUVjqBKXZw2tNuE5YceG = 1'b1; i2IIQfdSjOGJ0HAlaZdYe = 1'b0; end end 2'b10 : begin xSW8arCNXsyV5zIEXuGUQB = 2'b10; t69iUVjqBKXZw2tNuE5YceG = 1'b1; if (m0Pt9awzMYrRUb1BRHcMLqG) begin if (JomiEQo6ylRrlhLJPFsQTG == 1'b1) begin xSW8arCNXsyV5zIEXuGUQB = 2'b00; t69iUVjqBKXZw2tNuE5YceG = 1'b0; i2IIQfdSjOGJ0HAlaZdYe = 1'b0; end else begin i2IIQfdSjOGJ0HAlaZdYe = 1'b1; end end end default : begin xSW8arCNXsyV5zIEXuGUQB = 2'b00; i2IIQfdSjOGJ0HAlaZdYe = 1'b0; t69iUVjqBKXZw2tNuE5YceG = 1'b0; end endcase euwYuFBjOyzJ1StMM7x9lB = GP01IUV0xObQQCSdqL463C; qhMTHhfDKHqjrVnmTgdY6 = pDYTWTp6fyrEdA1XnDiP6E; pBYDq5TsLLci7qFUEEbLfB = Xf88wK4mkniJ6qfkmOXy2C; end assign g1oJwDFAtNAcPvLahTlMEB = euwYuFBjOyzJ1StMM7x9lB; assign wf5f4XnltnQYt1bEDWEp0F = n40UqkH7P32znVloyhHzXD; assign Q7D2KKVRLkwEPktPhyCkSD = qhMTHhfDKHqjrVnmTgdY6; endmodule