`timescale 1 ns / 1 ns module kkELk45BoVareqHanLSiwD (rstb, v04pHKxyc2sPW047bbyUgE, vLtlRIKgN8j1pwmLLNsPG, JzMAX1dysSuDOcRjDKM6jE, mFPagULjpfgerkfoXcLj6E, ZxXeSJVdqJaLdxkVQHDcKE, m5wgqFuUcW1FOMsh4Ru6H, KMtac8skVU06MkqFCILXMF, n3sKmw6MRNFgYu3FVurx4gF, ruH3uKgP1LYhGZv6tkbvYB, h5UJTRfxlrAz6m3sECIknXE, Fr5Lz9pdsoRhxTCNFip6AE, uG1VLsSqDTRiixegby6clE, qqi4ViVQH4ZOVdWVypt4yB, UKo8akspo4h0jsZ6g712NB, zzBKVZ6VX4ht5u9x9EjCiD, j83GXtGY1eMU252JJ6B9mC, r7Q5mFJeRMLiOPMHQDcQQB, wtshVXYU5akP8bsJW8meZH, w2g8aZ7DNLiB7xd9ema9tID, EpypH5ZIz8rvw2qkajrEUD, k5yT5mPpUVKMKN3fkRm1LR, hfxEgMPHtdNs5za4aJfZR); input rstb; input v04pHKxyc2sPW047bbyUgE; input [16:0] vLtlRIKgN8j1pwmLLNsPG; input [16:0] JzMAX1dysSuDOcRjDKM6jE; input [16:0] mFPagULjpfgerkfoXcLj6E; input [16:0] ZxXeSJVdqJaLdxkVQHDcKE; input signed [15:0] m5wgqFuUcW1FOMsh4Ru6H; input signed [15:0] KMtac8skVU06MkqFCILXMF; input signed [15:0] n3sKmw6MRNFgYu3FVurx4gF; input signed [15:0] ruH3uKgP1LYhGZv6tkbvYB; input signed [15:0] h5UJTRfxlrAz6m3sECIknXE; input signed [15:0] Fr5Lz9pdsoRhxTCNFip6AE; input signed [15:0] uG1VLsSqDTRiixegby6clE; input signed [15:0] qqi4ViVQH4ZOVdWVypt4yB; input UKo8akspo4h0jsZ6g712NB; output signed [15:0] zzBKVZ6VX4ht5u9x9EjCiD; output signed [15:0] j83GXtGY1eMU252JJ6B9mC; output signed [15:0] r7Q5mFJeRMLiOPMHQDcQQB; output signed [15:0] wtshVXYU5akP8bsJW8meZH; output signed [15:0] w2g8aZ7DNLiB7xd9ema9tID; output signed [15:0] EpypH5ZIz8rvw2qkajrEUD; output signed [15:0] k5yT5mPpUVKMKN3fkRm1LR; output signed [15:0] hfxEgMPHtdNs5za4aJfZR; wire signed [15:0] wQtS2qaE78f3Y1DG1Pi2cE; wire signed [15:0] TSiEK9Y9LFP93eIwf9K32F; wire signed [15:0] qqYA02t5VUHMdvk0DbMiIH; wire signed [15:0] vBlMyrCgC22Fut5ut8eC5F; wire signed [15:0] FfFNZ9spFyXrNhrofDq67G; wire signed [15:0] gTB5A1alvjs1wgYYkqPav; wire signed [15:0] YapR4aqvLec1XwDmzqE9KH; wire signed [15:0] W0accAMrUD2AeFMHHvYsF; wire fPxWcS5Nys1WvBWSYWvJrG; zVydWOLm2SZCpbjeNcZUmCpp #(.AddrWidth(17), .DataWidth(16) ) E7biabxSLcPGNoKkmdQk6C (.rstb(rstb), .v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .QDJhCuX1glwonJutj0sIMH(m5wgqFuUcW1FOMsh4Ru6H), .g0hVqHZpe6H7t41TOVwtoTE(h5UJTRfxlrAz6m3sECIknXE), .qmEenX2Yt9VTzGvbielz5B(vLtlRIKgN8j1pwmLLNsPG), .DiF2KV4VbJn3P66sh0MYvH(UKo8akspo4h0jsZ6g712NB), .ds3UaO1QhyfiWT7RZKX23G(wQtS2qaE78f3Y1DG1Pi2cE), .tCCvu1nsVn6k0oKnEbNi9E(TSiEK9Y9LFP93eIwf9K32F) ); assign zzBKVZ6VX4ht5u9x9EjCiD = wQtS2qaE78f3Y1DG1Pi2cE; zVydWOLm2SZCpbjeNcZUmCpp #(.AddrWidth(17), .DataWidth(16) ) oJl3TH6gWe25fGMscW3Da (.rstb(rstb), .v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .QDJhCuX1glwonJutj0sIMH(KMtac8skVU06MkqFCILXMF), .g0hVqHZpe6H7t41TOVwtoTE(Fr5Lz9pdsoRhxTCNFip6AE), .qmEenX2Yt9VTzGvbielz5B(JzMAX1dysSuDOcRjDKM6jE), .DiF2KV4VbJn3P66sh0MYvH(UKo8akspo4h0jsZ6g712NB), .ds3UaO1QhyfiWT7RZKX23G(qqYA02t5VUHMdvk0DbMiIH), .tCCvu1nsVn6k0oKnEbNi9E(vBlMyrCgC22Fut5ut8eC5F) ); assign j83GXtGY1eMU252JJ6B9mC = qqYA02t5VUHMdvk0DbMiIH; zVydWOLm2SZCpbjeNcZUmCpp #(.AddrWidth(17), .DataWidth(16) ) R4BJmTEufmjpXWftkSi9tG (.rstb(rstb), .v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .QDJhCuX1glwonJutj0sIMH(n3sKmw6MRNFgYu3FVurx4gF), .g0hVqHZpe6H7t41TOVwtoTE(uG1VLsSqDTRiixegby6clE), .qmEenX2Yt9VTzGvbielz5B(mFPagULjpfgerkfoXcLj6E), .DiF2KV4VbJn3P66sh0MYvH(UKo8akspo4h0jsZ6g712NB), .ds3UaO1QhyfiWT7RZKX23G(FfFNZ9spFyXrNhrofDq67G), .tCCvu1nsVn6k0oKnEbNi9E(gTB5A1alvjs1wgYYkqPav) ); assign r7Q5mFJeRMLiOPMHQDcQQB = FfFNZ9spFyXrNhrofDq67G; zVydWOLm2SZCpbjeNcZUmCpp #(.AddrWidth(17), .DataWidth(16) ) NyG7YBTWRpTZHuoR9Wtr5E (.rstb(rstb), .v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .QDJhCuX1glwonJutj0sIMH(ruH3uKgP1LYhGZv6tkbvYB), .g0hVqHZpe6H7t41TOVwtoTE(qqi4ViVQH4ZOVdWVypt4yB), .qmEenX2Yt9VTzGvbielz5B(ZxXeSJVdqJaLdxkVQHDcKE), .DiF2KV4VbJn3P66sh0MYvH(UKo8akspo4h0jsZ6g712NB), .ds3UaO1QhyfiWT7RZKX23G(YapR4aqvLec1XwDmzqE9KH), .tCCvu1nsVn6k0oKnEbNi9E(W0accAMrUD2AeFMHHvYsF) ); assign wtshVXYU5akP8bsJW8meZH = YapR4aqvLec1XwDmzqE9KH; assign w2g8aZ7DNLiB7xd9ema9tID = TSiEK9Y9LFP93eIwf9K32F; assign EpypH5ZIz8rvw2qkajrEUD = vBlMyrCgC22Fut5ut8eC5F; assign k5yT5mPpUVKMKN3fkRm1LR = gTB5A1alvjs1wgYYkqPav; assign hfxEgMPHtdNs5za4aJfZR = W0accAMrUD2AeFMHHvYsF; endmodule
