`timescale 1 ns / 1 ns module e61uBMMOD8obk5m2QBgMSL (v04pHKxyc2sPW047bbyUgE, JAMOfrNHxGSYDF0urqkLN, c070CKvbOwMMYffRzNpxjuG, pLZcRyd2lMVX3oSoEEblZE, R6zf5iqRNVEGVBO8egq8kF, BZMbpSF4BAilhRWeHczrfC, Ax88y9n8GnrKjg0yG0FKzE, CosmSfOlF9hl7OPB7KnKvB, rFrTP2XEQaUmbjytbnblxB); input v04pHKxyc2sPW047bbyUgE; input JAMOfrNHxGSYDF0urqkLN; input c070CKvbOwMMYffRzNpxjuG; input pLZcRyd2lMVX3oSoEEblZE; input R6zf5iqRNVEGVBO8egq8kF; output [5:0] BZMbpSF4BAilhRWeHczrfC; output Ax88y9n8GnrKjg0yG0FKzE; output CosmSfOlF9hl7OPB7KnKvB; output rFrTP2XEQaUmbjytbnblxB; reg [5:0] JomiEQo6ylRrlhLJPFsQTG; reg [1:0] X7FJ0jgk6hqdMN8BingGvE; reg [1:0] WXS42gmgDxS46057b3AGD; reg [5:0] GP01IUV0xObQQCSdqL463C; reg pDYTWTp6fyrEdA1XnDiP6E; reg [1:0] mb13NdjIe7rpJDLNih8AaE; reg Xf88wK4mkniJ6qfkmOXy2C; reg [5:0] i2IIQfdSjOGJ0HAlaZdYe; reg [1:0] xSW8arCNXsyV5zIEXuGUQB; reg [1:0] ck9Ya76HU61qWvvl3qwfRG; reg [5:0] dQhJtS5aSGZCPWaJqkkHi; reg t69iUVjqBKXZw2tNuE5YceG; reg [1:0] BNI9VucWF1TWsCAM4sBCHE; reg EIfu64RX7LMQGnynQeCGuD; reg [5:0] WX7lHFo8W3ZpxbqMsSFGGH; reg nNTCt2rbPOMpxZJonUxJrF; reg C24ghXBbSmP5ZsWcoJv4iD; reg XeR1BLGhFsA5XvRQUnMKDB; wire UZ4UUnX6yzJl5Maerfk2yC; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : h6oTzWU1a3otHwaiji95ID if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin JomiEQo6ylRrlhLJPFsQTG <= 6'b000000; GP01IUV0xObQQCSdqL463C <= 6'b000000; X7FJ0jgk6hqdMN8BingGvE <= 2'b00; WXS42gmgDxS46057b3AGD <= 2'b00; mb13NdjIe7rpJDLNih8AaE <= 2'b00; pDYTWTp6fyrEdA1XnDiP6E <= 1'b0; Xf88wK4mkniJ6qfkmOXy2C <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin JomiEQo6ylRrlhLJPFsQTG <= 6'b000000; GP01IUV0xObQQCSdqL463C <= 6'b000000; X7FJ0jgk6hqdMN8BingGvE <= 2'b00; WXS42gmgDxS46057b3AGD <= 2'b00; mb13NdjIe7rpJDLNih8AaE <= 2'b00; pDYTWTp6fyrEdA1XnDiP6E <= 1'b0; Xf88wK4mkniJ6qfkmOXy2C <= 1'b0; end else begin JomiEQo6ylRrlhLJPFsQTG <= i2IIQfdSjOGJ0HAlaZdYe; X7FJ0jgk6hqdMN8BingGvE <= xSW8arCNXsyV5zIEXuGUQB; WXS42gmgDxS46057b3AGD <= ck9Ya76HU61qWvvl3qwfRG; GP01IUV0xObQQCSdqL463C <= dQhJtS5aSGZCPWaJqkkHi; pDYTWTp6fyrEdA1XnDiP6E <= t69iUVjqBKXZw2tNuE5YceG; mb13NdjIe7rpJDLNih8AaE <= BNI9VucWF1TWsCAM4sBCHE; Xf88wK4mkniJ6qfkmOXy2C <= EIfu64RX7LMQGnynQeCGuD; end end end always @(GP01IUV0xObQQCSdqL463C, JomiEQo6ylRrlhLJPFsQTG, WXS42gmgDxS46057b3AGD, X7FJ0jgk6hqdMN8BingGvE, Xf88wK4mkniJ6qfkmOXy2C, c070CKvbOwMMYffRzNpxjuG, mb13NdjIe7rpJDLNih8AaE, pDYTWTp6fyrEdA1XnDiP6E, pLZcRyd2lMVX3oSoEEblZE) begin i2IIQfdSjOGJ0HAlaZdYe = JomiEQo6ylRrlhLJPFsQTG; xSW8arCNXsyV5zIEXuGUQB = X7FJ0jgk6hqdMN8BingGvE; ck9Ya76HU61qWvvl3qwfRG = WXS42gmgDxS46057b3AGD; dQhJtS5aSGZCPWaJqkkHi = GP01IUV0xObQQCSdqL463C; t69iUVjqBKXZw2tNuE5YceG = pDYTWTp6fyrEdA1XnDiP6E; BNI9VucWF1TWsCAM4sBCHE = mb13NdjIe7rpJDLNih8AaE; EIfu64RX7LMQGnynQeCGuD = Xf88wK4mkniJ6qfkmOXy2C; case ( mb13NdjIe7rpJDLNih8AaE) 2'b00 : begin BNI9VucWF1TWsCAM4sBCHE = 2'b00; EIfu64RX7LMQGnynQeCGuD = 1'b0; if (WXS42gmgDxS46057b3AGD == 2'b01) begin BNI9VucWF1TWsCAM4sBCHE = 2'b01; end end 2'b01 : begin EIfu64RX7LMQGnynQeCGuD = 1'b0; if (WXS42gmgDxS46057b3AGD == 2'b10) begin BNI9VucWF1TWsCAM4sBCHE = 2'b10; end end 2'b10 : begin EIfu64RX7LMQGnynQeCGuD = 1'b0; if (WXS42gmgDxS46057b3AGD == 2'b01) begin BNI9VucWF1TWsCAM4sBCHE = 2'b11; EIfu64RX7LMQGnynQeCGuD = 1'b1; end end 2'b11 : begin if (WXS42gmgDxS46057b3AGD == 2'b01) begin BNI9VucWF1TWsCAM4sBCHE = 2'b11; EIfu64RX7LMQGnynQeCGuD = 1'b1; end else begin EIfu64RX7LMQGnynQeCGuD = 1'b0; BNI9VucWF1TWsCAM4sBCHE = 2'b00; end end default : begin BNI9VucWF1TWsCAM4sBCHE = 2'b00; EIfu64RX7LMQGnynQeCGuD = 1'b0; end endcase case ( WXS42gmgDxS46057b3AGD) 2'b00 : begin ck9Ya76HU61qWvvl3qwfRG = 2'b00; dQhJtS5aSGZCPWaJqkkHi = 6'b000000; nNTCt2rbPOMpxZJonUxJrF = 1'b0; if (c070CKvbOwMMYffRzNpxjuG && (JomiEQo6ylRrlhLJPFsQTG == 6'b111111)) begin ck9Ya76HU61qWvvl3qwfRG = 2'b01; end end 2'b01 : begin ck9Ya76HU61qWvvl3qwfRG = 2'b01; nNTCt2rbPOMpxZJonUxJrF = pLZcRyd2lMVX3oSoEEblZE; if (pLZcRyd2lMVX3oSoEEblZE) begin if (GP01IUV0xObQQCSdqL463C == 6'b111111) begin ck9Ya76HU61qWvvl3qwfRG = 2'b10; end dQhJtS5aSGZCPWaJqkkHi = GP01IUV0xObQQCSdqL463C + 6'b000001; end end 2'b10 : begin nNTCt2rbPOMpxZJonUxJrF = 1'b1; if (GP01IUV0xObQQCSdqL463C == 6'b111111) begin if (c070CKvbOwMMYffRzNpxjuG && (JomiEQo6ylRrlhLJPFsQTG == 6'b111111)) begin ck9Ya76HU61qWvvl3qwfRG = 2'b01; end else begin ck9Ya76HU61qWvvl3qwfRG = 2'b00; end end dQhJtS5aSGZCPWaJqkkHi = GP01IUV0xObQQCSdqL463C + 6'b000001; end default : begin ck9Ya76HU61qWvvl3qwfRG = 2'b00; dQhJtS5aSGZCPWaJqkkHi = 6'b000000; nNTCt2rbPOMpxZJonUxJrF = 1'b0; end endcase case ( X7FJ0jgk6hqdMN8BingGvE) 2'b00 : begin xSW8arCNXsyV5zIEXuGUQB = 2'b00; i2IIQfdSjOGJ0HAlaZdYe = 6'b000000; t69iUVjqBKXZw2tNuE5YceG = 1'b0; if (c070CKvbOwMMYffRzNpxjuG) begin xSW8arCNXsyV5zIEXuGUQB = 2'b01; i2IIQfdSjOGJ0HAlaZdYe = 6'b000001; end end 2'b01 : begin xSW8arCNXsyV5zIEXuGUQB = 2'b01; t69iUVjqBKXZw2tNuE5YceG = 1'b0; if (c070CKvbOwMMYffRzNpxjuG) begin if (JomiEQo6ylRrlhLJPFsQTG == 6'b111111) begin xSW8arCNXsyV5zIEXuGUQB = 2'b10; t69iUVjqBKXZw2tNuE5YceG = 1'b1; end else begin xSW8arCNXsyV5zIEXuGUQB = 2'b01; end i2IIQfdSjOGJ0HAlaZdYe = JomiEQo6ylRrlhLJPFsQTG + 6'b000001; end end 2'b10 : begin xSW8arCNXsyV5zIEXuGUQB = 2'b10; if (c070CKvbOwMMYffRzNpxjuG) begin if (JomiEQo6ylRrlhLJPFsQTG == 6'b111111) begin xSW8arCNXsyV5zIEXuGUQB = 2'b01; t69iUVjqBKXZw2tNuE5YceG = 1'b0; end else begin xSW8arCNXsyV5zIEXuGUQB = 2'b10; t69iUVjqBKXZw2tNuE5YceG = 1'b1; end i2IIQfdSjOGJ0HAlaZdYe = JomiEQo6ylRrlhLJPFsQTG + 6'b000001; end end default : begin xSW8arCNXsyV5zIEXuGUQB = 2'b00; i2IIQfdSjOGJ0HAlaZdYe = 6'b111111; t69iUVjqBKXZw2tNuE5YceG = 1'b0; end endcase WX7lHFo8W3ZpxbqMsSFGGH = GP01IUV0xObQQCSdqL463C; C24ghXBbSmP5ZsWcoJv4iD = pDYTWTp6fyrEdA1XnDiP6E; XeR1BLGhFsA5XvRQUnMKDB = Xf88wK4mkniJ6qfkmOXy2C; end assign BZMbpSF4BAilhRWeHczrfC = WX7lHFo8W3ZpxbqMsSFGGH; assign Ax88y9n8GnrKjg0yG0FKzE = nNTCt2rbPOMpxZJonUxJrF; assign CosmSfOlF9hl7OPB7KnKvB = C24ghXBbSmP5ZsWcoJv4iD; assign rFrTP2XEQaUmbjytbnblxB = XeR1BLGhFsA5XvRQUnMKDB; endmodule