`timescale 1 ns / 1 ns module c5frKpr1OF9l0qPiwsMhI2 (v04pHKxyc2sPW047bbyUgE, JAMOfrNHxGSYDF0urqkLN, kIsHJAwQMWbIiCsXfX1rTG, DKGIysOp4cb2Wy4ifYHB8D, R6zf5iqRNVEGVBO8egq8kF, yTf5WZbZOLm2uKwJmXk5sG, wGlnEfCkRPxniOjCaZH6XG, RDvlVEJspE7WkJvNmR8a6C); input v04pHKxyc2sPW047bbyUgE; input JAMOfrNHxGSYDF0urqkLN; input kIsHJAwQMWbIiCsXfX1rTG; input DKGIysOp4cb2Wy4ifYHB8D; input R6zf5iqRNVEGVBO8egq8kF; output yTf5WZbZOLm2uKwJmXk5sG; output wGlnEfCkRPxniOjCaZH6XG; output RDvlVEJspE7WkJvNmR8a6C; reg [1:0] X7FJ0jgk6hqdMN8BingGvE; reg [1:0] WXS42gmgDxS46057b3AGD; reg GP01IUV0xObQQCSdqL463C; reg [1:0] mb13NdjIe7rpJDLNih8AaE; reg [1:0] xSW8arCNXsyV5zIEXuGUQB; reg [1:0] ck9Ya76HU61qWvvl3qwfRG; reg dQhJtS5aSGZCPWaJqkkHi; reg [1:0] BNI9VucWF1TWsCAM4sBCHE; reg f0LoJaVTftOyaXbKcYjRST; reg udLm1gCfK1bsBCzyYOebLD; reg mjQQDV7qVUmtyjMgSHu2bC; reg S86yDRz3lzvCeFmkKizFJD; wire vYr9oPWf1tgVRPgCssDAtD; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : h6oTzWU1a3otHwaiji95ID if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin GP01IUV0xObQQCSdqL463C <= 1'b0; X7FJ0jgk6hqdMN8BingGvE <= 2'b00; WXS42gmgDxS46057b3AGD <= 2'b00; mb13NdjIe7rpJDLNih8AaE <= 2'b00; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin GP01IUV0xObQQCSdqL463C <= 1'b0; X7FJ0jgk6hqdMN8BingGvE <= 2'b00; WXS42gmgDxS46057b3AGD <= 2'b00; mb13NdjIe7rpJDLNih8AaE <= 2'b00; end else begin X7FJ0jgk6hqdMN8BingGvE <= xSW8arCNXsyV5zIEXuGUQB; WXS42gmgDxS46057b3AGD <= ck9Ya76HU61qWvvl3qwfRG; GP01IUV0xObQQCSdqL463C <= dQhJtS5aSGZCPWaJqkkHi; mb13NdjIe7rpJDLNih8AaE <= BNI9VucWF1TWsCAM4sBCHE; end end end always @(DKGIysOp4cb2Wy4ifYHB8D, GP01IUV0xObQQCSdqL463C, WXS42gmgDxS46057b3AGD, X7FJ0jgk6hqdMN8BingGvE, kIsHJAwQMWbIiCsXfX1rTG, mb13NdjIe7rpJDLNih8AaE) begin xSW8arCNXsyV5zIEXuGUQB = X7FJ0jgk6hqdMN8BingGvE; ck9Ya76HU61qWvvl3qwfRG = WXS42gmgDxS46057b3AGD; dQhJtS5aSGZCPWaJqkkHi = GP01IUV0xObQQCSdqL463C; BNI9VucWF1TWsCAM4sBCHE = mb13NdjIe7rpJDLNih8AaE; case ( mb13NdjIe7rpJDLNih8AaE) 2'b00 : begin BNI9VucWF1TWsCAM4sBCHE = 2'b00; S86yDRz3lzvCeFmkKizFJD = 1'b0; if (WXS42gmgDxS46057b3AGD == 2'b01) begin BNI9VucWF1TWsCAM4sBCHE = 2'b01; end end 2'b01 : begin S86yDRz3lzvCeFmkKizFJD = 1'b0; if (WXS42gmgDxS46057b3AGD == 2'b00) begin BNI9VucWF1TWsCAM4sBCHE = 2'b10; end end 2'b10 : begin S86yDRz3lzvCeFmkKizFJD = 1'b0; if ((X7FJ0jgk6hqdMN8BingGvE == 2'b11) && kIsHJAwQMWbIiCsXfX1rTG) begin BNI9VucWF1TWsCAM4sBCHE = 2'b11; end end 2'b11 : begin S86yDRz3lzvCeFmkKizFJD = 1'b1; if (DKGIysOp4cb2Wy4ifYHB8D) begin BNI9VucWF1TWsCAM4sBCHE = 2'b00; end end default : begin BNI9VucWF1TWsCAM4sBCHE = 2'b00; S86yDRz3lzvCeFmkKizFJD = 1'b0; end endcase case ( WXS42gmgDxS46057b3AGD) 2'b00 : begin ck9Ya76HU61qWvvl3qwfRG = 2'b00; dQhJtS5aSGZCPWaJqkkHi = 1'b0; udLm1gCfK1bsBCzyYOebLD = 1'b0; if ((X7FJ0jgk6hqdMN8BingGvE == 2'b11) && kIsHJAwQMWbIiCsXfX1rTG) begin ck9Ya76HU61qWvvl3qwfRG = 2'b01; udLm1gCfK1bsBCzyYOebLD = DKGIysOp4cb2Wy4ifYHB8D; end end 2'b01 : begin udLm1gCfK1bsBCzyYOebLD = DKGIysOp4cb2Wy4ifYHB8D; if (DKGIysOp4cb2Wy4ifYHB8D) begin ck9Ya76HU61qWvvl3qwfRG = 2'b00; end end default : begin ck9Ya76HU61qWvvl3qwfRG = 2'b00; dQhJtS5aSGZCPWaJqkkHi = 1'b0; udLm1gCfK1bsBCzyYOebLD = 1'b0; end endcase case ( X7FJ0jgk6hqdMN8BingGvE) 2'b00 : begin xSW8arCNXsyV5zIEXuGUQB = 2'b00; mjQQDV7qVUmtyjMgSHu2bC = 1'b0; if (kIsHJAwQMWbIiCsXfX1rTG) begin xSW8arCNXsyV5zIEXuGUQB = 2'b11; end end 2'b11 : begin xSW8arCNXsyV5zIEXuGUQB = 2'b11; mjQQDV7qVUmtyjMgSHu2bC = 1'b0; if (kIsHJAwQMWbIiCsXfX1rTG) begin xSW8arCNXsyV5zIEXuGUQB = 2'b10; mjQQDV7qVUmtyjMgSHu2bC = 1'b1; end end 2'b10 : begin mjQQDV7qVUmtyjMgSHu2bC = 1'b0; xSW8arCNXsyV5zIEXuGUQB = 2'b10; if (kIsHJAwQMWbIiCsXfX1rTG) begin xSW8arCNXsyV5zIEXuGUQB = 2'b11; end end default : begin xSW8arCNXsyV5zIEXuGUQB = 2'b00; mjQQDV7qVUmtyjMgSHu2bC = 1'b0; end endcase f0LoJaVTftOyaXbKcYjRST = GP01IUV0xObQQCSdqL463C; end assign yTf5WZbZOLm2uKwJmXk5sG = f0LoJaVTftOyaXbKcYjRST; assign wGlnEfCkRPxniOjCaZH6XG = udLm1gCfK1bsBCzyYOebLD; assign RDvlVEJspE7WkJvNmR8a6C = mjQQDV7qVUmtyjMgSHu2bC; endmodule