`timescale 1 ns / 1 ns module m0wR0p8t3oV06dM5Osycg9 (v04pHKxyc2sPW047bbyUgE, JAMOfrNHxGSYDF0urqkLN, DZol1WsbVnSldsei0SiI9E, sIaC8spfzCmUwexq8stmB, R6zf5iqRNVEGVBO8egq8kF, zqdZMmoxIs9zmnL4kATVuC, a8rK4qdEuNCWHLdYbR2f8, O6TgnxqnGk692qEmnZQFTC, XfCDnggI1Y1qaMzSOLL0TD); input v04pHKxyc2sPW047bbyUgE; input JAMOfrNHxGSYDF0urqkLN; input DZol1WsbVnSldsei0SiI9E; input sIaC8spfzCmUwexq8stmB; input R6zf5iqRNVEGVBO8egq8kF; output zqdZMmoxIs9zmnL4kATVuC; output a8rK4qdEuNCWHLdYbR2f8; output O6TgnxqnGk692qEmnZQFTC; output XfCDnggI1Y1qaMzSOLL0TD; reg JomiEQo6ylRrlhLJPFsQTG; reg [1:0] X7FJ0jgk6hqdMN8BingGvE; reg [1:0] WXS42gmgDxS46057b3AGD; reg GP01IUV0xObQQCSdqL463C; reg pDYTWTp6fyrEdA1XnDiP6E; reg [1:0] mb13NdjIe7rpJDLNih8AaE; reg Xf88wK4mkniJ6qfkmOXy2C; reg i2IIQfdSjOGJ0HAlaZdYe; reg [1:0] xSW8arCNXsyV5zIEXuGUQB; reg [1:0] ck9Ya76HU61qWvvl3qwfRG; reg dQhJtS5aSGZCPWaJqkkHi; reg t69iUVjqBKXZw2tNuE5YceG; reg [1:0] BNI9VucWF1TWsCAM4sBCHE; reg EIfu64RX7LMQGnynQeCGuD; reg FTmbjaPeOhErAS6D1MUlWB; reg gSX2i71vFz3rrbsDU0gsUF; reg pJQMR6eedLw0JCRx8qs1KE; reg f5wnPIXmY4DkSIOQfFS2MB; wire DXTyywsKoi0LpqWz2bUNwH; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : h6oTzWU1a3otHwaiji95ID if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin JomiEQo6ylRrlhLJPFsQTG <= 1'b0; GP01IUV0xObQQCSdqL463C <= 1'b0; X7FJ0jgk6hqdMN8BingGvE <= 2'b00; WXS42gmgDxS46057b3AGD <= 2'b00; mb13NdjIe7rpJDLNih8AaE <= 2'b00; pDYTWTp6fyrEdA1XnDiP6E <= 1'b0; Xf88wK4mkniJ6qfkmOXy2C <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin JomiEQo6ylRrlhLJPFsQTG <= 1'b0; GP01IUV0xObQQCSdqL463C <= 1'b0; X7FJ0jgk6hqdMN8BingGvE <= 2'b00; WXS42gmgDxS46057b3AGD <= 2'b00; mb13NdjIe7rpJDLNih8AaE <= 2'b00; pDYTWTp6fyrEdA1XnDiP6E <= 1'b0; Xf88wK4mkniJ6qfkmOXy2C <= 1'b0; end else begin JomiEQo6ylRrlhLJPFsQTG <= i2IIQfdSjOGJ0HAlaZdYe; X7FJ0jgk6hqdMN8BingGvE <= xSW8arCNXsyV5zIEXuGUQB; WXS42gmgDxS46057b3AGD <= ck9Ya76HU61qWvvl3qwfRG; GP01IUV0xObQQCSdqL463C <= dQhJtS5aSGZCPWaJqkkHi; pDYTWTp6fyrEdA1XnDiP6E <= t69iUVjqBKXZw2tNuE5YceG; mb13NdjIe7rpJDLNih8AaE <= BNI9VucWF1TWsCAM4sBCHE; Xf88wK4mkniJ6qfkmOXy2C <= EIfu64RX7LMQGnynQeCGuD; end end end always @(DZol1WsbVnSldsei0SiI9E, GP01IUV0xObQQCSdqL463C, JomiEQo6ylRrlhLJPFsQTG, WXS42gmgDxS46057b3AGD, X7FJ0jgk6hqdMN8BingGvE, Xf88wK4mkniJ6qfkmOXy2C, mb13NdjIe7rpJDLNih8AaE, pDYTWTp6fyrEdA1XnDiP6E, sIaC8spfzCmUwexq8stmB) begin i2IIQfdSjOGJ0HAlaZdYe = JomiEQo6ylRrlhLJPFsQTG; xSW8arCNXsyV5zIEXuGUQB = X7FJ0jgk6hqdMN8BingGvE; ck9Ya76HU61qWvvl3qwfRG = WXS42gmgDxS46057b3AGD; dQhJtS5aSGZCPWaJqkkHi = GP01IUV0xObQQCSdqL463C; t69iUVjqBKXZw2tNuE5YceG = pDYTWTp6fyrEdA1XnDiP6E; BNI9VucWF1TWsCAM4sBCHE = mb13NdjIe7rpJDLNih8AaE; EIfu64RX7LMQGnynQeCGuD = Xf88wK4mkniJ6qfkmOXy2C; case ( mb13NdjIe7rpJDLNih8AaE) 2'b00 : begin BNI9VucWF1TWsCAM4sBCHE = 2'b00; EIfu64RX7LMQGnynQeCGuD = 1'b0; if (WXS42gmgDxS46057b3AGD == 2'b01) begin BNI9VucWF1TWsCAM4sBCHE = 2'b01; end end 2'b01 : begin EIfu64RX7LMQGnynQeCGuD = ! (GP01IUV0xObQQCSdqL463C == 1'b0); if (WXS42gmgDxS46057b3AGD == 2'b10) begin BNI9VucWF1TWsCAM4sBCHE = 2'b10; end end 2'b10 : begin EIfu64RX7LMQGnynQeCGuD = 1'b0; if (WXS42gmgDxS46057b3AGD == 2'b01) begin BNI9VucWF1TWsCAM4sBCHE = 2'b11; end end 2'b11 : begin if (WXS42gmgDxS46057b3AGD == 2'b01) begin BNI9VucWF1TWsCAM4sBCHE = 2'b11; EIfu64RX7LMQGnynQeCGuD = ! (GP01IUV0xObQQCSdqL463C == 1'b0); end else begin EIfu64RX7LMQGnynQeCGuD = 1'b0; BNI9VucWF1TWsCAM4sBCHE = 2'b00; end end default : begin BNI9VucWF1TWsCAM4sBCHE = 2'b00; EIfu64RX7LMQGnynQeCGuD = 1'b0; end endcase case ( WXS42gmgDxS46057b3AGD) 2'b00 : begin ck9Ya76HU61qWvvl3qwfRG = 2'b00; dQhJtS5aSGZCPWaJqkkHi = 1'b0; gSX2i71vFz3rrbsDU0gsUF = 1'b0; if (pDYTWTp6fyrEdA1XnDiP6E) begin ck9Ya76HU61qWvvl3qwfRG = 2'b01; gSX2i71vFz3rrbsDU0gsUF = sIaC8spfzCmUwexq8stmB; if (sIaC8spfzCmUwexq8stmB) begin dQhJtS5aSGZCPWaJqkkHi = 1'b1; end end end 2'b01 : begin ck9Ya76HU61qWvvl3qwfRG = 2'b01; gSX2i71vFz3rrbsDU0gsUF = sIaC8spfzCmUwexq8stmB; if (sIaC8spfzCmUwexq8stmB) begin if (GP01IUV0xObQQCSdqL463C == 1'b1) begin ck9Ya76HU61qWvvl3qwfRG = 2'b10; dQhJtS5aSGZCPWaJqkkHi = 1'b0; end else begin dQhJtS5aSGZCPWaJqkkHi = 1'b1; end end end 2'b10 : begin gSX2i71vFz3rrbsDU0gsUF = 1'b0; if (GP01IUV0xObQQCSdqL463C == 1'b1) begin dQhJtS5aSGZCPWaJqkkHi = 1'b0; if (pDYTWTp6fyrEdA1XnDiP6E) begin ck9Ya76HU61qWvvl3qwfRG = 2'b01; end else begin ck9Ya76HU61qWvvl3qwfRG = 2'b00; end end else begin dQhJtS5aSGZCPWaJqkkHi = 1'b1; end end default : begin ck9Ya76HU61qWvvl3qwfRG = 2'b00; dQhJtS5aSGZCPWaJqkkHi = 1'b0; gSX2i71vFz3rrbsDU0gsUF = 1'b0; end endcase case ( X7FJ0jgk6hqdMN8BingGvE) 2'b00 : begin xSW8arCNXsyV5zIEXuGUQB = 2'b00; i2IIQfdSjOGJ0HAlaZdYe = 1'b0; t69iUVjqBKXZw2tNuE5YceG = 1'b0; if (DZol1WsbVnSldsei0SiI9E) begin xSW8arCNXsyV5zIEXuGUQB = 2'b01; i2IIQfdSjOGJ0HAlaZdYe = 1'b1; end end 2'b01 : begin xSW8arCNXsyV5zIEXuGUQB = 2'b01; t69iUVjqBKXZw2tNuE5YceG = 1'b0; if (DZol1WsbVnSldsei0SiI9E) begin xSW8arCNXsyV5zIEXuGUQB = 2'b10; t69iUVjqBKXZw2tNuE5YceG = 1'b1; i2IIQfdSjOGJ0HAlaZdYe = 1'b0; end end 2'b10 : begin xSW8arCNXsyV5zIEXuGUQB = 2'b10; t69iUVjqBKXZw2tNuE5YceG = 1'b1; if (DZol1WsbVnSldsei0SiI9E) begin if (JomiEQo6ylRrlhLJPFsQTG == 1'b1) begin xSW8arCNXsyV5zIEXuGUQB = 2'b00; t69iUVjqBKXZw2tNuE5YceG = 1'b0; i2IIQfdSjOGJ0HAlaZdYe = 1'b0; end else begin i2IIQfdSjOGJ0HAlaZdYe = 1'b1; end end end default : begin xSW8arCNXsyV5zIEXuGUQB = 2'b00; i2IIQfdSjOGJ0HAlaZdYe = 1'b0; t69iUVjqBKXZw2tNuE5YceG = 1'b0; end endcase FTmbjaPeOhErAS6D1MUlWB = GP01IUV0xObQQCSdqL463C; pJQMR6eedLw0JCRx8qs1KE = pDYTWTp6fyrEdA1XnDiP6E; f5wnPIXmY4DkSIOQfFS2MB = Xf88wK4mkniJ6qfkmOXy2C; end assign zqdZMmoxIs9zmnL4kATVuC = FTmbjaPeOhErAS6D1MUlWB; assign a8rK4qdEuNCWHLdYbR2f8 = gSX2i71vFz3rrbsDU0gsUF; assign O6TgnxqnGk692qEmnZQFTC = pJQMR6eedLw0JCRx8qs1KE; assign XfCDnggI1Y1qaMzSOLL0TD = f5wnPIXmY4DkSIOQfFS2MB; endmodule