`timescale 1 ns / 1 ns module yzoOoF7555t5sVm5WeZ9lC (v04pHKxyc2sPW047bbyUgE, JAMOfrNHxGSYDF0urqkLN, j8MMagsoA5t6IysA2ZD3X4F, k3VfrgkD6DWITJL9WW5W4D, pPn6MVGqBLqJ0xzN2WYfFG, OUMqBzkN19EDa2VTABMa2E, qbEnMIxMUsx8pYkF1gFd7D, jNZ4xylBKAANfCL11XNxzB, R6zf5iqRNVEGVBO8egq8kF, VWSiqDgxQN9a2J7zRy3p4E, LhqlKpPzANkuN2xC8HYciC, s1N0USypDrc4xyzxc4XEMr, sZ7bCwrhIAA80IOhzh695); input v04pHKxyc2sPW047bbyUgE; input JAMOfrNHxGSYDF0urqkLN; input j8MMagsoA5t6IysA2ZD3X4F; input signed [15:0] k3VfrgkD6DWITJL9WW5W4D; input signed [15:0] pPn6MVGqBLqJ0xzN2WYfFG; input signed [15:0] OUMqBzkN19EDa2VTABMa2E; input signed [15:0] qbEnMIxMUsx8pYkF1gFd7D; input jNZ4xylBKAANfCL11XNxzB; input R6zf5iqRNVEGVBO8egq8kF; output signed [15:0] VWSiqDgxQN9a2J7zRy3p4E; output signed [15:0] LhqlKpPzANkuN2xC8HYciC; output signed [15:0] s1N0USypDrc4xyzxc4XEMr; output signed [15:0] sZ7bCwrhIAA80IOhzh695; reg AxdzJminNkFCybtxxeC5hH; reg signed [16:0] p9Q1ZdD8IyrQGhwT1XXpAwH; reg signed [16:0] FrouE4YVttOqChzztq9MRG; reg signed [16:0] i4FJCC6Xft9yUijVwpyTC0E; reg signed [16:0] N5RqGyuQKrj2dkBK5NIpfD; reg b8PGIsG3FsdAJqb7hOUD1oC; reg signed [16:0] u6qmTF9ijEkH9xmDrm95pEF; reg signed [16:0] MP4qvH0uMShcprYVFxKkUD; reg signed [16:0] COyf11G22yt2ahr9Ucug2E; reg signed [16:0] bYOlGODgGA4hK2uJ9g4xaG; reg signed [15:0] aydyoHsGbz0wVGlm34qlsB; reg signed [15:0] H0BpAwmwCivCDsbLQ5qvCC; reg signed [15:0] aRq4LmGEDdp6eFXcSQc6HE; reg signed [15:0] WZvcQ1OGi1O0JWI4mdwqx; reg Pq4nKEqqr18aLXK1kX1dfH; reg signed [16:0] a6WUK3shR7OoXJD6OQBcnbC; reg signed [16:0] z8sdLNMywEyzxM9eSpPklMB; reg signed [16:0] x4JZ8sOjxjZWNeN08B95t5B; reg signed [16:0] JpNj7HaVF5ISgAz8d6xCmE; reg signed [16:0] lyJA6GgUdA5yMT3KGmkiBB; reg signed [16:0] YTn6r1K2cbi4BzelKHgZMH; reg signed [16:0] T6fhnGgnCx4gzNMLRlfJsB; reg signed [16:0] QaUWOROgNo7uvlOzzIL7gF; reg signed [16:0] f9uiVizQ8iG3TggFQMEaqMB; reg signed [16:0] whyOPXTaiRJEg5hgsaLJCG; reg signed [16:0] yqGXdE6pHXRFGlXkfvbpKC; reg signed [16:0] UzOnWFVNmsGSUzlrKfHqwF; reg signed [16:0] b9p1O84anZ1REVMvdH9T6cE; reg signed [16:0] uOyZcxygSH2ObqTFvmjZLD; reg signed [16:0] giifcHhQs1eZ2W9VasanfG; reg signed [16:0] Ht14IixEv7IQddUNB8FBaF; reg signed [16:0] g64FBA6XTYfJB3gQdH04OJH; reg signed [16:0] cefQ41MlYs7FI4dPMnads; reg signed [16:0] ZLjCoy1mhX7nS8r36AkTnG; reg signed [16:0] z6qazKI7KMGAFLe2KGVVFE; reg signed [16:0] xE4ft4QLMQrp1NtpcdoU2D; reg signed [16:0] b3b6q6yOnUzkdBZha4J35NB; reg signed [16:0] xsDfZ2jarysSjALlotRtW; reg signed [16:0] YLWHYhSBwDrFHhQzmw106G; reg signed [16:0] J3I5o2R6c9ixHmw1Oa9EvE; reg signed [16:0] bN7pv94LbbUjIRAxJt4lf; reg signed [16:0] PZRWIojv1r4p0mRa5bnL8G; reg signed [16:0] iZxjhcD6M6J4jJWVBLDvjG; wire PbKVjWnrIoG3VeFj7j32fF; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : aMdxH72OgWBZw20gQc6DxE if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin AxdzJminNkFCybtxxeC5hH <= 1'b0; p9Q1ZdD8IyrQGhwT1XXpAwH <= 17'sb00000000000000000; FrouE4YVttOqChzztq9MRG <= 17'sb00000000000000000; i4FJCC6Xft9yUijVwpyTC0E <= 17'sb00000000000000000; N5RqGyuQKrj2dkBK5NIpfD <= 17'sb00000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin AxdzJminNkFCybtxxeC5hH <= 1'b0; p9Q1ZdD8IyrQGhwT1XXpAwH <= 17'sb00000000000000000; FrouE4YVttOqChzztq9MRG <= 17'sb00000000000000000; i4FJCC6Xft9yUijVwpyTC0E <= 17'sb00000000000000000; N5RqGyuQKrj2dkBK5NIpfD <= 17'sb00000000000000000; end else begin AxdzJminNkFCybtxxeC5hH <= b8PGIsG3FsdAJqb7hOUD1oC; p9Q1ZdD8IyrQGhwT1XXpAwH <= u6qmTF9ijEkH9xmDrm95pEF; FrouE4YVttOqChzztq9MRG <= MP4qvH0uMShcprYVFxKkUD; i4FJCC6Xft9yUijVwpyTC0E <= COyf11G22yt2ahr9Ucug2E; N5RqGyuQKrj2dkBK5NIpfD <= bYOlGODgGA4hK2uJ9g4xaG; end end end always @(AxdzJminNkFCybtxxeC5hH, FrouE4YVttOqChzztq9MRG, N5RqGyuQKrj2dkBK5NIpfD, OUMqBzkN19EDa2VTABMa2E, i4FJCC6Xft9yUijVwpyTC0E, j8MMagsoA5t6IysA2ZD3X4F, jNZ4xylBKAANfCL11XNxzB, k3VfrgkD6DWITJL9WW5W4D, p9Q1ZdD8IyrQGhwT1XXpAwH, pPn6MVGqBLqJ0xzN2WYfFG, qbEnMIxMUsx8pYkF1gFd7D) begin b9p1O84anZ1REVMvdH9T6cE = 17'sb00000000000000000; uOyZcxygSH2ObqTFvmjZLD = 17'sb00000000000000000; giifcHhQs1eZ2W9VasanfG = 17'sb00000000000000000; Ht14IixEv7IQddUNB8FBaF = 17'sb00000000000000000; g64FBA6XTYfJB3gQdH04OJH = 17'sb00000000000000000; cefQ41MlYs7FI4dPMnads = 17'sb00000000000000000; ZLjCoy1mhX7nS8r36AkTnG = 17'sb00000000000000000; z6qazKI7KMGAFLe2KGVVFE = 17'sb00000000000000000; xE4ft4QLMQrp1NtpcdoU2D = 17'sb00000000000000000; b3b6q6yOnUzkdBZha4J35NB = 17'sb00000000000000000; xsDfZ2jarysSjALlotRtW = 17'sb00000000000000000; YLWHYhSBwDrFHhQzmw106G = 17'sb00000000000000000; J3I5o2R6c9ixHmw1Oa9EvE = 17'sb00000000000000000; bN7pv94LbbUjIRAxJt4lf = 17'sb00000000000000000; PZRWIojv1r4p0mRa5bnL8G = 17'sb00000000000000000; iZxjhcD6M6J4jJWVBLDvjG = 17'sb00000000000000000; u6qmTF9ijEkH9xmDrm95pEF = p9Q1ZdD8IyrQGhwT1XXpAwH; MP4qvH0uMShcprYVFxKkUD = FrouE4YVttOqChzztq9MRG; COyf11G22yt2ahr9Ucug2E = i4FJCC6Xft9yUijVwpyTC0E; bYOlGODgGA4hK2uJ9g4xaG = N5RqGyuQKrj2dkBK5NIpfD; b8PGIsG3FsdAJqb7hOUD1oC = jNZ4xylBKAANfCL11XNxzB; if (j8MMagsoA5t6IysA2ZD3X4F != 1'b0) begin if (jNZ4xylBKAANfCL11XNxzB) begin b9p1O84anZ1REVMvdH9T6cE = {k3VfrgkD6DWITJL9WW5W4D[15], k3VfrgkD6DWITJL9WW5W4D}; uOyZcxygSH2ObqTFvmjZLD = {qbEnMIxMUsx8pYkF1gFd7D[15], qbEnMIxMUsx8pYkF1gFd7D}; u6qmTF9ijEkH9xmDrm95pEF = b9p1O84anZ1REVMvdH9T6cE + uOyZcxygSH2ObqTFvmjZLD; giifcHhQs1eZ2W9VasanfG = {k3VfrgkD6DWITJL9WW5W4D[15], k3VfrgkD6DWITJL9WW5W4D}; Ht14IixEv7IQddUNB8FBaF = {qbEnMIxMUsx8pYkF1gFd7D[15], qbEnMIxMUsx8pYkF1gFd7D}; COyf11G22yt2ahr9Ucug2E = giifcHhQs1eZ2W9VasanfG - Ht14IixEv7IQddUNB8FBaF; g64FBA6XTYfJB3gQdH04OJH = {pPn6MVGqBLqJ0xzN2WYfFG[15], pPn6MVGqBLqJ0xzN2WYfFG}; cefQ41MlYs7FI4dPMnads = {OUMqBzkN19EDa2VTABMa2E[15], OUMqBzkN19EDa2VTABMa2E}; bYOlGODgGA4hK2uJ9g4xaG = g64FBA6XTYfJB3gQdH04OJH + cefQ41MlYs7FI4dPMnads; ZLjCoy1mhX7nS8r36AkTnG = {pPn6MVGqBLqJ0xzN2WYfFG[15], pPn6MVGqBLqJ0xzN2WYfFG}; z6qazKI7KMGAFLe2KGVVFE = {OUMqBzkN19EDa2VTABMa2E[15], OUMqBzkN19EDa2VTABMa2E}; MP4qvH0uMShcprYVFxKkUD = ZLjCoy1mhX7nS8r36AkTnG - z6qazKI7KMGAFLe2KGVVFE; end end else if (jNZ4xylBKAANfCL11XNxzB) begin xE4ft4QLMQrp1NtpcdoU2D = {k3VfrgkD6DWITJL9WW5W4D[15], k3VfrgkD6DWITJL9WW5W4D}; b3b6q6yOnUzkdBZha4J35NB = {OUMqBzkN19EDa2VTABMa2E[15], OUMqBzkN19EDa2VTABMa2E}; u6qmTF9ijEkH9xmDrm95pEF = xE4ft4QLMQrp1NtpcdoU2D + b3b6q6yOnUzkdBZha4J35NB; xsDfZ2jarysSjALlotRtW = {k3VfrgkD6DWITJL9WW5W4D[15], k3VfrgkD6DWITJL9WW5W4D}; YLWHYhSBwDrFHhQzmw106G = {OUMqBzkN19EDa2VTABMa2E[15], OUMqBzkN19EDa2VTABMa2E}; COyf11G22yt2ahr9Ucug2E = xsDfZ2jarysSjALlotRtW - YLWHYhSBwDrFHhQzmw106G; J3I5o2R6c9ixHmw1Oa9EvE = {pPn6MVGqBLqJ0xzN2WYfFG[15], pPn6MVGqBLqJ0xzN2WYfFG}; bN7pv94LbbUjIRAxJt4lf = {qbEnMIxMUsx8pYkF1gFd7D[15], qbEnMIxMUsx8pYkF1gFd7D}; MP4qvH0uMShcprYVFxKkUD = J3I5o2R6c9ixHmw1Oa9EvE + bN7pv94LbbUjIRAxJt4lf; PZRWIojv1r4p0mRa5bnL8G = {pPn6MVGqBLqJ0xzN2WYfFG[15], pPn6MVGqBLqJ0xzN2WYfFG}; iZxjhcD6M6J4jJWVBLDvjG = {qbEnMIxMUsx8pYkF1gFd7D[15], qbEnMIxMUsx8pYkF1gFd7D}; bYOlGODgGA4hK2uJ9g4xaG = PZRWIojv1r4p0mRa5bnL8G - iZxjhcD6M6J4jJWVBLDvjG; end a6WUK3shR7OoXJD6OQBcnbC = ({p9Q1ZdD8IyrQGhwT1XXpAwH[16], p9Q1ZdD8IyrQGhwT1XXpAwH[16:1]}) + $signed({1'b0, p9Q1ZdD8IyrQGhwT1XXpAwH[0]}); z8sdLNMywEyzxM9eSpPklMB = a6WUK3shR7OoXJD6OQBcnbC >>> 8'd1; x4JZ8sOjxjZWNeN08B95t5B = {z8sdLNMywEyzxM9eSpPklMB[15:0], 1'b0}; aydyoHsGbz0wVGlm34qlsB = x4JZ8sOjxjZWNeN08B95t5B[15:0]; JpNj7HaVF5ISgAz8d6xCmE = ({FrouE4YVttOqChzztq9MRG[16], FrouE4YVttOqChzztq9MRG[16:1]}) + $signed({1'b0, FrouE4YVttOqChzztq9MRG[0]}); lyJA6GgUdA5yMT3KGmkiBB = JpNj7HaVF5ISgAz8d6xCmE >>> 8'd1; YTn6r1K2cbi4BzelKHgZMH = {lyJA6GgUdA5yMT3KGmkiBB[15:0], 1'b0}; H0BpAwmwCivCDsbLQ5qvCC = YTn6r1K2cbi4BzelKHgZMH[15:0]; T6fhnGgnCx4gzNMLRlfJsB = ({i4FJCC6Xft9yUijVwpyTC0E[16], i4FJCC6Xft9yUijVwpyTC0E[16:1]}) + $signed({1'b0, i4FJCC6Xft9yUijVwpyTC0E[0]}); QaUWOROgNo7uvlOzzIL7gF = T6fhnGgnCx4gzNMLRlfJsB >>> 8'd1; f9uiVizQ8iG3TggFQMEaqMB = {QaUWOROgNo7uvlOzzIL7gF[15:0], 1'b0}; aRq4LmGEDdp6eFXcSQc6HE = f9uiVizQ8iG3TggFQMEaqMB[15:0]; whyOPXTaiRJEg5hgsaLJCG = ({N5RqGyuQKrj2dkBK5NIpfD[16], N5RqGyuQKrj2dkBK5NIpfD[16:1]}) + $signed({1'b0, N5RqGyuQKrj2dkBK5NIpfD[0]}); yqGXdE6pHXRFGlXkfvbpKC = whyOPXTaiRJEg5hgsaLJCG >>> 8'd1; UzOnWFVNmsGSUzlrKfHqwF = {yqGXdE6pHXRFGlXkfvbpKC[15:0], 1'b0}; WZvcQ1OGi1O0JWI4mdwqx = UzOnWFVNmsGSUzlrKfHqwF[15:0]; Pq4nKEqqr18aLXK1kX1dfH = AxdzJminNkFCybtxxeC5hH; end assign VWSiqDgxQN9a2J7zRy3p4E = aydyoHsGbz0wVGlm34qlsB; assign LhqlKpPzANkuN2xC8HYciC = H0BpAwmwCivCDsbLQ5qvCC; assign s1N0USypDrc4xyzxc4XEMr = aRq4LmGEDdp6eFXcSQc6HE; assign sZ7bCwrhIAA80IOhzh695 = WZvcQ1OGi1O0JWI4mdwqx; endmodule