`timescale 1 ns / 1 ns module bLNpla6dKRnNqV9xT7W46B (v04pHKxyc2sPW047bbyUgE, JAMOfrNHxGSYDF0urqkLN, S6Ue4SxCiz8dBHTO2guOUE, POhLmCr6emegQDte8TzyQ, E9kfQ0vBTIumIk9ATubhJH, GFkF4uUefeRBOH9Wes3V5D, NdNevEoWljk83nSbsGDU1C, Tf0EDmJTni9HuTSAYQFT2F, qp9pmnimi6dV0X7tI2Wt6B, Gw5sPQAOzFLVF06eF1AOGF, uO7PvkjtbrbcoMU62rs5JF, R6zf5iqRNVEGVBO8egq8kF, qmhLAZZAHFrO09l1zXnPRC, JMtgCMT5TVzyJSn9uILA1, xYJCS7zMCKI1yYR3Bx1XrD, AaqUpSvCGAV1YR86nIsLWH); input v04pHKxyc2sPW047bbyUgE; input JAMOfrNHxGSYDF0urqkLN; input signed [15:0] S6Ue4SxCiz8dBHTO2guOUE; input signed [15:0] POhLmCr6emegQDte8TzyQ; input signed [15:0] E9kfQ0vBTIumIk9ATubhJH; input signed [15:0] GFkF4uUefeRBOH9Wes3V5D; input NdNevEoWljk83nSbsGDU1C; input signed [15:0] Tf0EDmJTni9HuTSAYQFT2F; input signed [15:0] qp9pmnimi6dV0X7tI2Wt6B; input signed [15:0] Gw5sPQAOzFLVF06eF1AOGF; input signed [15:0] uO7PvkjtbrbcoMU62rs5JF; input R6zf5iqRNVEGVBO8egq8kF; output signed [15:0] qmhLAZZAHFrO09l1zXnPRC; output signed [15:0] JMtgCMT5TVzyJSn9uILA1; output signed [15:0] xYJCS7zMCKI1yYR3Bx1XrD; output signed [15:0] AaqUpSvCGAV1YR86nIsLWH; reg signed [15:0] XOQBCWZyBA9fPc87mG5IsD; reg signed [15:0] jgpSuUOXE6beAUY2P4Iv4C; reg signed [15:0] s6mgKiePlUcVLouID5veYH; reg signed [15:0] W3WuRCFnI5ngJZRPIZcluH; reg signed [15:0] PJ83Ne7TovKBk1QalAPkbF; reg signed [15:0] PQB4vyiY2hzUb277RaVY2G; reg mBEavkbBsOgXvycfTD0hMD; reg mRiDGTkFKo4RMA0LJKgthG; reg KmAm4o6cjyOTvVGRHZ5CwE; reg signed [15:0] Y4G0Jzpc0pu9WjWBN3cG3G; reg signed [15:0] yi5TBCH5TW5biX3U7QsRqE; reg signed [15:0] UV2a0iFkGBexVZbqWWEZtH; reg signed [15:0] srmdhX8C2dssNj53K6bvXB; reg signed [15:0] PI4X2832OFOysxpHuBiM9G; reg signed [15:0] wBO6oB2d6g6Z4IwDoFEshF; reg JRIoLUeCq9mXSVlgE57gFE; reg tSpBSFRas5hrgrmHKg0BzD; reg SNSO4dX03KiNOAsJChroeG; wire lEeKsyOAQXjFKEeD6pbdWF; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : MczQYJ6MT1pYZD7C1UhQv if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin XOQBCWZyBA9fPc87mG5IsD <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin XOQBCWZyBA9fPc87mG5IsD <= 16'sb0000000000000000; end else begin XOQBCWZyBA9fPc87mG5IsD <= S6Ue4SxCiz8dBHTO2guOUE; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : xwyxj2YIc64Lxvl4r8S8mG if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin jgpSuUOXE6beAUY2P4Iv4C <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin jgpSuUOXE6beAUY2P4Iv4C <= 16'sb0000000000000000; end else begin jgpSuUOXE6beAUY2P4Iv4C <= XOQBCWZyBA9fPc87mG5IsD; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : L1HBH8O5DRbGBa9XvBX70C if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin s6mgKiePlUcVLouID5veYH <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin s6mgKiePlUcVLouID5veYH <= 16'sb0000000000000000; end else begin s6mgKiePlUcVLouID5veYH <= jgpSuUOXE6beAUY2P4Iv4C; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : s2CWr6rrksK4W7N0omU97HD if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin W3WuRCFnI5ngJZRPIZcluH <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin W3WuRCFnI5ngJZRPIZcluH <= 16'sb0000000000000000; end else begin W3WuRCFnI5ngJZRPIZcluH <= POhLmCr6emegQDte8TzyQ; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : k1Zsi6BUVrSUjLbIYwh26G if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin PJ83Ne7TovKBk1QalAPkbF <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin PJ83Ne7TovKBk1QalAPkbF <= 16'sb0000000000000000; end else begin PJ83Ne7TovKBk1QalAPkbF <= W3WuRCFnI5ngJZRPIZcluH; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : TPi3Fu9uFLztbkFwa0H53D if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin PQB4vyiY2hzUb277RaVY2G <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin PQB4vyiY2hzUb277RaVY2G <= 16'sb0000000000000000; end else begin PQB4vyiY2hzUb277RaVY2G <= PJ83Ne7TovKBk1QalAPkbF; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : IBmSJmjQmOQZECy1AykU1D if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin mBEavkbBsOgXvycfTD0hMD <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin mBEavkbBsOgXvycfTD0hMD <= 1'b0; end else begin mBEavkbBsOgXvycfTD0hMD <= NdNevEoWljk83nSbsGDU1C; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : VNPcEW4KZxpAtEz0DCT8vD if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin mRiDGTkFKo4RMA0LJKgthG <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin mRiDGTkFKo4RMA0LJKgthG <= 1'b0; end else begin mRiDGTkFKo4RMA0LJKgthG <= mBEavkbBsOgXvycfTD0hMD; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : t8uWAeIAh3IMbN9UNxoYBKD if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin KmAm4o6cjyOTvVGRHZ5CwE <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin KmAm4o6cjyOTvVGRHZ5CwE <= 1'b0; end else begin KmAm4o6cjyOTvVGRHZ5CwE <= mRiDGTkFKo4RMA0LJKgthG; end end end BalZ6iNPh05BZIILLQfca k6VwTDKyQk0wkkUi6c3ojtC (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .s6mgKiePlUcVLouID5veYH(s6mgKiePlUcVLouID5veYH), .PQB4vyiY2hzUb277RaVY2G(PQB4vyiY2hzUb277RaVY2G), .KmAm4o6cjyOTvVGRHZ5CwE(KmAm4o6cjyOTvVGRHZ5CwE), .Tf0EDmJTni9HuTSAYQFT2F(Tf0EDmJTni9HuTSAYQFT2F), .qp9pmnimi6dV0X7tI2Wt6B(qp9pmnimi6dV0X7tI2Wt6B), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .qmhLAZZAHFrO09l1zXnPRC(qmhLAZZAHFrO09l1zXnPRC), .JMtgCMT5TVzyJSn9uILA1(JMtgCMT5TVzyJSn9uILA1) ); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : QtzxgwI206U33aXvIkKdwD if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin Y4G0Jzpc0pu9WjWBN3cG3G <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin Y4G0Jzpc0pu9WjWBN3cG3G <= 16'sb0000000000000000; end else begin Y4G0Jzpc0pu9WjWBN3cG3G <= E9kfQ0vBTIumIk9ATubhJH; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : awX33YTQEl2OxkV2HHm04D if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin yi5TBCH5TW5biX3U7QsRqE <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin yi5TBCH5TW5biX3U7QsRqE <= 16'sb0000000000000000; end else begin yi5TBCH5TW5biX3U7QsRqE <= Y4G0Jzpc0pu9WjWBN3cG3G; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : wroVmvZXsLz1H55Ur0PrpB if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin UV2a0iFkGBexVZbqWWEZtH <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin UV2a0iFkGBexVZbqWWEZtH <= 16'sb0000000000000000; end else begin UV2a0iFkGBexVZbqWWEZtH <= yi5TBCH5TW5biX3U7QsRqE; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : z8NMcVNSFzdoHNpSsC5DBLF if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin srmdhX8C2dssNj53K6bvXB <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin srmdhX8C2dssNj53K6bvXB <= 16'sb0000000000000000; end else begin srmdhX8C2dssNj53K6bvXB <= GFkF4uUefeRBOH9Wes3V5D; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : j2gHN9roTaQcXLtCUWIL9F if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin PI4X2832OFOysxpHuBiM9G <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin PI4X2832OFOysxpHuBiM9G <= 16'sb0000000000000000; end else begin PI4X2832OFOysxpHuBiM9G <= srmdhX8C2dssNj53K6bvXB; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : eVDXDpbSTruDFXBM6ygPaB if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin wBO6oB2d6g6Z4IwDoFEshF <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin wBO6oB2d6g6Z4IwDoFEshF <= 16'sb0000000000000000; end else begin wBO6oB2d6g6Z4IwDoFEshF <= PI4X2832OFOysxpHuBiM9G; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : a2bprYW6bhaVvTUhwUfmVQF if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin JRIoLUeCq9mXSVlgE57gFE <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin JRIoLUeCq9mXSVlgE57gFE <= 1'b0; end else begin JRIoLUeCq9mXSVlgE57gFE <= NdNevEoWljk83nSbsGDU1C; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : RfFhiu7TcZArCuQWZZoVsB if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin tSpBSFRas5hrgrmHKg0BzD <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin tSpBSFRas5hrgrmHKg0BzD <= 1'b0; end else begin tSpBSFRas5hrgrmHKg0BzD <= JRIoLUeCq9mXSVlgE57gFE; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : owLoaMKUokO7uUwJJovpJE if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin SNSO4dX03KiNOAsJChroeG <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin SNSO4dX03KiNOAsJChroeG <= 1'b0; end else begin SNSO4dX03KiNOAsJChroeG <= tSpBSFRas5hrgrmHKg0BzD; end end end wD13SKguCvt6FPikYT4rmB JOQQNSibUv7LmaKv3pf63F (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .UV2a0iFkGBexVZbqWWEZtH(UV2a0iFkGBexVZbqWWEZtH), .wBO6oB2d6g6Z4IwDoFEshF(wBO6oB2d6g6Z4IwDoFEshF), .SNSO4dX03KiNOAsJChroeG(SNSO4dX03KiNOAsJChroeG), .Gw5sPQAOzFLVF06eF1AOGF(Gw5sPQAOzFLVF06eF1AOGF), .uO7PvkjtbrbcoMU62rs5JF(uO7PvkjtbrbcoMU62rs5JF), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .xYJCS7zMCKI1yYR3Bx1XrD(xYJCS7zMCKI1yYR3Bx1XrD), .AaqUpSvCGAV1YR86nIsLWH(AaqUpSvCGAV1YR86nIsLWH) ); endmodule