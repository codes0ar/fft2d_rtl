`timescale 1 ns / 1 ns module LB48BKt395PB3Xbcuwg3wC (v04pHKxyc2sPW047bbyUgE, JAMOfrNHxGSYDF0urqkLN, DbYwoM2JCYD9mwcRRKmb6G, WbySmFpEqdJe6nrpd6KgG, pCWATI9lTIGbmXTtLuLAGB, yTf5WZbZOLm2uKwJmXk5sG, wGlnEfCkRPxniOjCaZH6XG, i4y6Td18s9Zr0JbepLQtjC, k3FlrGNoOUOhUgHDIDYGouE, RDvlVEJspE7WkJvNmR8a6C, R6zf5iqRNVEGVBO8egq8kF, t30W3eeadZl9O9RnQCafyED, flGpcmOyc38fKmqiV5eQvF); input v04pHKxyc2sPW047bbyUgE; input JAMOfrNHxGSYDF0urqkLN; input signed [15:0] DbYwoM2JCYD9mwcRRKmb6G; input signed [15:0] WbySmFpEqdJe6nrpd6KgG; input pCWATI9lTIGbmXTtLuLAGB; input yTf5WZbZOLm2uKwJmXk5sG; input wGlnEfCkRPxniOjCaZH6XG; input signed [15:0] i4y6Td18s9Zr0JbepLQtjC; input signed [15:0] k3FlrGNoOUOhUgHDIDYGouE; input RDvlVEJspE7WkJvNmR8a6C; input R6zf5iqRNVEGVBO8egq8kF; output signed [15:0] t30W3eeadZl9O9RnQCafyED; output signed [15:0] flGpcmOyc38fKmqiV5eQvF; wire signed [15:0] x3T5ivGGBQbBK8kZOoMj3; wire signed [15:0] cMIOWiDVVCoNgM2IifcBEE; wire j4o2xcEQspSUTgY2fvzdEdD; reg de21duRLbf27relCAO1YZB; wire signed [15:0] N2ZdE4zLlq5uRV4rcE2wdE; wire signed [15:0] iOhy3XYM3su7ndksftfCZG; wire AECH0r3KnKo0RJFepDhYUD; wire twcuYIJzeZMBjyHmZ1FZDD; reg signed [15:0] jCeVBfgGpg4ODtaTTQIgZH; reg signed [15:0] lI5eRWU0Hmm71ItlHz1XD; reg signed [15:0] p8q8wLTlQG0dlPaw6UilCB; reg signed [15:0] CxgFTw1cIpgtTBm0G0iIGE; reg signed [15:0] hZ6V0Vos1jyuJExMLN1ea; reg signed [15:0] TzSfIMdbsYlfcbdYVDW7IE; reg signed [15:0] XMU8TKFj7fRDeSlFsaP4eC; reg signed [15:0] wU64i77CqFqKfsCs2glSxC; reg signed [15:0] nBWi8KlMIOvUV5djMbF0CD; reg signed [15:0] m0RTEXqA15w9eP2jMaxNBoD; reg signed [15:0] OvRzP6mVEGIsekLbBoFXkF; reg signed [15:0] zd5MqAnK6OPkumgkpYCpQF; reg signed [15:0] csMK1iTp18g0vZYjmk9JZD; reg signed [15:0] dTkGd8OUQ83dmglc4Bt8vF; reg signed [16:0] wFsaSfYltg6TlrWqY1FyGE; reg signed [16:0] T5BRwctOUS2khp8Rzx4l9; reg signed [16:0] t1ZySna7c411biAKwiSaOlF; reg signed [16:0] d8074IV5GByVrE9OuVeZYRF; reg signed [15:0] f6eYgeW0rCfd0LIvc2SGHB; reg signed [15:0] m5VNx3xnw67GgdN5661tXkG; reg signed [15:0] IMsvh2kSL36ZxgH6ovKFz; reg signed [15:0] ZvsdK7IB0VkAxGNAOwtzgD; reg q6XydGshj15r9Fju4CQ2iT; reg KuSB40UBeOqvdWcrRv76OB; wire signed [16:0] kHkm1dHei7pqznzynbBKwE; wire signed [16:0] Oym0ZQxbxCKFQ5X3kAuPi; wire signed [16:0] YIMNIvC4K9LQaGT0TCHkcE; wire signed [16:0] IQG3jvRoS6AY8QAkGyV9b; wire signed [16:0] g4G8R7TlPZ9NvGqBSUmdb7F; wire signed [16:0] ndTxZ4yEyGpSsXjLwP10HB; wire signed [16:0] plZaC1IiHJbFqqHndxJpKC; wire signed [16:0] B8fYUIF4y2YvoVPCpuCb0; wire signed [16:0] Yb4qpWQhiQpsJ5laLdw1dG; wire signed [16:0] XETUnhSmrTZNec4mfH5bhE; wire signed [16:0] krcDen5cyZ3crTZ2yfXap; wire signed [16:0] fpzEAgYwqhsLsJYv4qlk8E; wire signed [16:0] n0J4kP9YDHfDkhTNLn56dJ; wire signed [16:0] UpDw6anZs0bMPETxgXld9F; wire signed [16:0] b31KhkrKeVwOtEcPIkvs3; wire signed [16:0] Lcbc8UkQ7CVMIZTyIGqp7G; wire signed [16:0] KinlMSwCRgZdG2BmpRDJAG; wire signed [16:0] t1uTFhJAosQhy0vBWGPplXD; wire signed [16:0] Pr2dhfiX07pLlRUhRGiSR; wire signed [16:0] LgvxMrXuJRlmlCyhLVJYyE; wire signed [16:0] ATjS2KECQ0ZiH7CL8LEnE; wire signed [16:0] RPKurxOe2f65XPpdjKRZMF; wire signed [16:0] a2Lel9XzXgLNrkI13pSAHKE; wire signed [16:0] VJAT39ZYYYO4RWA7Qqf56F; reg signed [15:0] mgknRxAcgFrHqTt5CZvnSF; reg signed [15:0] sCFM4WicR6deeSAdSwumP; reg BKNY6GzA6oGZumjzTATycD; wire signed [15:0] uUcj3UAzjmPW47yNyzbT8C; wire signed [15:0] uwZv0qzQLi0MDBWLWzKuAG; wire n65LdbEr6NMNaEFcjX8Fh6F; wire signed [15:0] x9j7a5gok64zzNKnvdJNnE; wire signed [15:0] bPL0FcLvoxhO0amTUOV9QC; wire signed [15:0] r4JngA0ZVhEElGRZci9fohF; wire signed [15:0] a8xx20Fc5nKc8DbqSwNBuB; reg vLT6ef7BJliTDpt4k5jqF; wire nePc9BiseLZlqhuLXpwEvG; r0u9EENf7w7dFzlB1BYZL7F ftPsaxEa6Qv5RNEVVRTJoH (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .DbYwoM2JCYD9mwcRRKmb6G(DbYwoM2JCYD9mwcRRKmb6G), .WbySmFpEqdJe6nrpd6KgG(WbySmFpEqdJe6nrpd6KgG), .pCWATI9lTIGbmXTtLuLAGB(pCWATI9lTIGbmXTtLuLAGB), .i4y6Td18s9Zr0JbepLQtjC(i4y6Td18s9Zr0JbepLQtjC), .k3FlrGNoOUOhUgHDIDYGouE(k3FlrGNoOUOhUgHDIDYGouE), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .x3T5ivGGBQbBK8kZOoMj3(x3T5ivGGBQbBK8kZOoMj3), .cMIOWiDVVCoNgM2IifcBEE(cMIOWiDVVCoNgM2IifcBEE), .j4o2xcEQspSUTgY2fvzdEdD(j4o2xcEQspSUTgY2fvzdEdD) ); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : MczQYJ6MT1pYZD7C1UhQv if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin de21duRLbf27relCAO1YZB <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin de21duRLbf27relCAO1YZB <= 1'b0; end else begin de21duRLbf27relCAO1YZB <= wGlnEfCkRPxniOjCaZH6XG; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : ad105sTzL9xAsBGc6tDsQD if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin jCeVBfgGpg4ODtaTTQIgZH <= 16'sb0000000000000000; lI5eRWU0Hmm71ItlHz1XD <= 16'sb0000000000000000; p8q8wLTlQG0dlPaw6UilCB <= 16'sb0000000000000000; CxgFTw1cIpgtTBm0G0iIGE <= 16'sb0000000000000000; hZ6V0Vos1jyuJExMLN1ea <= 16'sb0000000000000000; TzSfIMdbsYlfcbdYVDW7IE <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin jCeVBfgGpg4ODtaTTQIgZH <= 16'sb0000000000000000; lI5eRWU0Hmm71ItlHz1XD <= 16'sb0000000000000000; p8q8wLTlQG0dlPaw6UilCB <= 16'sb0000000000000000; CxgFTw1cIpgtTBm0G0iIGE <= 16'sb0000000000000000; hZ6V0Vos1jyuJExMLN1ea <= 16'sb0000000000000000; TzSfIMdbsYlfcbdYVDW7IE <= 16'sb0000000000000000; end else begin jCeVBfgGpg4ODtaTTQIgZH <= XMU8TKFj7fRDeSlFsaP4eC; lI5eRWU0Hmm71ItlHz1XD <= wU64i77CqFqKfsCs2glSxC; p8q8wLTlQG0dlPaw6UilCB <= nBWi8KlMIOvUV5djMbF0CD; CxgFTw1cIpgtTBm0G0iIGE <= m0RTEXqA15w9eP2jMaxNBoD; hZ6V0Vos1jyuJExMLN1ea <= OvRzP6mVEGIsekLbBoFXkF; TzSfIMdbsYlfcbdYVDW7IE <= zd5MqAnK6OPkumgkpYCpQF; end end end always @(AECH0r3KnKo0RJFepDhYUD, CxgFTw1cIpgtTBm0G0iIGE, N2ZdE4zLlq5uRV4rcE2wdE, TzSfIMdbsYlfcbdYVDW7IE, hZ6V0Vos1jyuJExMLN1ea, iOhy3XYM3su7ndksftfCZG, jCeVBfgGpg4ODtaTTQIgZH, lI5eRWU0Hmm71ItlHz1XD, p8q8wLTlQG0dlPaw6UilCB, twcuYIJzeZMBjyHmZ1FZDD, yTf5WZbZOLm2uKwJmXk5sG) begin XMU8TKFj7fRDeSlFsaP4eC = jCeVBfgGpg4ODtaTTQIgZH; wU64i77CqFqKfsCs2glSxC = lI5eRWU0Hmm71ItlHz1XD; nBWi8KlMIOvUV5djMbF0CD = p8q8wLTlQG0dlPaw6UilCB; m0RTEXqA15w9eP2jMaxNBoD = CxgFTw1cIpgtTBm0G0iIGE; OvRzP6mVEGIsekLbBoFXkF = hZ6V0Vos1jyuJExMLN1ea; zd5MqAnK6OPkumgkpYCpQF = TzSfIMdbsYlfcbdYVDW7IE; if (yTf5WZbZOLm2uKwJmXk5sG) begin OvRzP6mVEGIsekLbBoFXkF = p8q8wLTlQG0dlPaw6UilCB; zd5MqAnK6OPkumgkpYCpQF = CxgFTw1cIpgtTBm0G0iIGE; end else begin OvRzP6mVEGIsekLbBoFXkF = jCeVBfgGpg4ODtaTTQIgZH; zd5MqAnK6OPkumgkpYCpQF = lI5eRWU0Hmm71ItlHz1XD; end if (twcuYIJzeZMBjyHmZ1FZDD) begin if (AECH0r3KnKo0RJFepDhYUD == 1'b1) begin nBWi8KlMIOvUV5djMbF0CD = N2ZdE4zLlq5uRV4rcE2wdE; m0RTEXqA15w9eP2jMaxNBoD = iOhy3XYM3su7ndksftfCZG; end else begin XMU8TKFj7fRDeSlFsaP4eC = N2ZdE4zLlq5uRV4rcE2wdE; wU64i77CqFqKfsCs2glSxC = iOhy3XYM3su7ndksftfCZG; end end csMK1iTp18g0vZYjmk9JZD = hZ6V0Vos1jyuJExMLN1ea; dTkGd8OUQ83dmglc4Bt8vF = TzSfIMdbsYlfcbdYVDW7IE; end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : plVzUyM9ssc0g5eFRKR67 if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin wFsaSfYltg6TlrWqY1FyGE <= 17'sb00000000000000000; T5BRwctOUS2khp8Rzx4l9 <= 17'sb00000000000000000; t1ZySna7c411biAKwiSaOlF <= 17'sb00000000000000000; d8074IV5GByVrE9OuVeZYRF <= 17'sb00000000000000000; mgknRxAcgFrHqTt5CZvnSF <= 16'sb0000000000000000; sCFM4WicR6deeSAdSwumP <= 16'sb0000000000000000; BKNY6GzA6oGZumjzTATycD <= 1'b0; f6eYgeW0rCfd0LIvc2SGHB <= 16'sb0000000000000000; m5VNx3xnw67GgdN5661tXkG <= 16'sb0000000000000000; IMsvh2kSL36ZxgH6ovKFz <= 16'sb0000000000000000; ZvsdK7IB0VkAxGNAOwtzgD <= 16'sb0000000000000000; q6XydGshj15r9Fju4CQ2iT <= 1'b0; KuSB40UBeOqvdWcrRv76OB <= 1'b0; vLT6ef7BJliTDpt4k5jqF <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin wFsaSfYltg6TlrWqY1FyGE <= 17'sb00000000000000000; T5BRwctOUS2khp8Rzx4l9 <= 17'sb00000000000000000; t1ZySna7c411biAKwiSaOlF <= 17'sb00000000000000000; d8074IV5GByVrE9OuVeZYRF <= 17'sb00000000000000000; mgknRxAcgFrHqTt5CZvnSF <= 16'sb0000000000000000; sCFM4WicR6deeSAdSwumP <= 16'sb0000000000000000; BKNY6GzA6oGZumjzTATycD <= 1'b0; f6eYgeW0rCfd0LIvc2SGHB <= 16'sb0000000000000000; m5VNx3xnw67GgdN5661tXkG <= 16'sb0000000000000000; IMsvh2kSL36ZxgH6ovKFz <= 16'sb0000000000000000; ZvsdK7IB0VkAxGNAOwtzgD <= 16'sb0000000000000000; q6XydGshj15r9Fju4CQ2iT <= 1'b0; KuSB40UBeOqvdWcrRv76OB <= 1'b0; vLT6ef7BJliTDpt4k5jqF <= 1'b0; end else begin wFsaSfYltg6TlrWqY1FyGE <= kHkm1dHei7pqznzynbBKwE; T5BRwctOUS2khp8Rzx4l9 <= Oym0ZQxbxCKFQ5X3kAuPi; t1ZySna7c411biAKwiSaOlF <= YIMNIvC4K9LQaGT0TCHkcE; d8074IV5GByVrE9OuVeZYRF <= IQG3jvRoS6AY8QAkGyV9b; vLT6ef7BJliTDpt4k5jqF <= KuSB40UBeOqvdWcrRv76OB; KuSB40UBeOqvdWcrRv76OB <= q6XydGshj15r9Fju4CQ2iT; IMsvh2kSL36ZxgH6ovKFz <= f6eYgeW0rCfd0LIvc2SGHB; ZvsdK7IB0VkAxGNAOwtzgD <= m5VNx3xnw67GgdN5661tXkG; f6eYgeW0rCfd0LIvc2SGHB <= x3T5ivGGBQbBK8kZOoMj3; m5VNx3xnw67GgdN5661tXkG <= cMIOWiDVVCoNgM2IifcBEE; mgknRxAcgFrHqTt5CZvnSF <= csMK1iTp18g0vZYjmk9JZD; sCFM4WicR6deeSAdSwumP <= dTkGd8OUQ83dmglc4Bt8vF; BKNY6GzA6oGZumjzTATycD <= de21duRLbf27relCAO1YZB; q6XydGshj15r9Fju4CQ2iT <= RDvlVEJspE7WkJvNmR8a6C && j4o2xcEQspSUTgY2fvzdEdD; end end end assign n65LdbEr6NMNaEFcjX8Fh6F = ( ! RDvlVEJspE7WkJvNmR8a6C) && j4o2xcEQspSUTgY2fvzdEdD; assign KinlMSwCRgZdG2BmpRDJAG = {csMK1iTp18g0vZYjmk9JZD[15], csMK1iTp18g0vZYjmk9JZD}; assign t1uTFhJAosQhy0vBWGPplXD = {IMsvh2kSL36ZxgH6ovKFz[15], IMsvh2kSL36ZxgH6ovKFz}; assign kHkm1dHei7pqznzynbBKwE = KinlMSwCRgZdG2BmpRDJAG + t1uTFhJAosQhy0vBWGPplXD; assign Pr2dhfiX07pLlRUhRGiSR = {csMK1iTp18g0vZYjmk9JZD[15], csMK1iTp18g0vZYjmk9JZD}; assign LgvxMrXuJRlmlCyhLVJYyE = {IMsvh2kSL36ZxgH6ovKFz[15], IMsvh2kSL36ZxgH6ovKFz}; assign YIMNIvC4K9LQaGT0TCHkcE = Pr2dhfiX07pLlRUhRGiSR - LgvxMrXuJRlmlCyhLVJYyE; assign ATjS2KECQ0ZiH7CL8LEnE = {dTkGd8OUQ83dmglc4Bt8vF[15], dTkGd8OUQ83dmglc4Bt8vF}; assign RPKurxOe2f65XPpdjKRZMF = {ZvsdK7IB0VkAxGNAOwtzgD[15], ZvsdK7IB0VkAxGNAOwtzgD}; assign Oym0ZQxbxCKFQ5X3kAuPi = ATjS2KECQ0ZiH7CL8LEnE + RPKurxOe2f65XPpdjKRZMF; assign a2Lel9XzXgLNrkI13pSAHKE = {dTkGd8OUQ83dmglc4Bt8vF[15], dTkGd8OUQ83dmglc4Bt8vF}; assign VJAT39ZYYYO4RWA7Qqf56F = {ZvsdK7IB0VkAxGNAOwtzgD[15], ZvsdK7IB0VkAxGNAOwtzgD}; assign IQG3jvRoS6AY8QAkGyV9b = a2Lel9XzXgLNrkI13pSAHKE - VJAT39ZYYYO4RWA7Qqf56F; assign uUcj3UAzjmPW47yNyzbT8C = x3T5ivGGBQbBK8kZOoMj3; assign uwZv0qzQLi0MDBWLWzKuAG = cMIOWiDVVCoNgM2IifcBEE; assign g4G8R7TlPZ9NvGqBSUmdb7F = ({wFsaSfYltg6TlrWqY1FyGE[16], wFsaSfYltg6TlrWqY1FyGE[16:1]}) + $signed({1'b0, wFsaSfYltg6TlrWqY1FyGE[0]}); assign ndTxZ4yEyGpSsXjLwP10HB = g4G8R7TlPZ9NvGqBSUmdb7F >>> 8'd1; assign plZaC1IiHJbFqqHndxJpKC = {ndTxZ4yEyGpSsXjLwP10HB[15:0], 1'b0}; assign x9j7a5gok64zzNKnvdJNnE = plZaC1IiHJbFqqHndxJpKC[15:0]; assign B8fYUIF4y2YvoVPCpuCb0 = ({T5BRwctOUS2khp8Rzx4l9[16], T5BRwctOUS2khp8Rzx4l9[16:1]}) + $signed({1'b0, T5BRwctOUS2khp8Rzx4l9[0]}); assign Yb4qpWQhiQpsJ5laLdw1dG = B8fYUIF4y2YvoVPCpuCb0 >>> 8'd1; assign XETUnhSmrTZNec4mfH5bhE = {Yb4qpWQhiQpsJ5laLdw1dG[15:0], 1'b0}; assign bPL0FcLvoxhO0amTUOV9QC = XETUnhSmrTZNec4mfH5bhE[15:0]; assign krcDen5cyZ3crTZ2yfXap = ({t1ZySna7c411biAKwiSaOlF[16], t1ZySna7c411biAKwiSaOlF[16:1]}) + $signed({1'b0, t1ZySna7c411biAKwiSaOlF[0]}); assign fpzEAgYwqhsLsJYv4qlk8E = krcDen5cyZ3crTZ2yfXap >>> 8'd1; assign n0J4kP9YDHfDkhTNLn56dJ = {fpzEAgYwqhsLsJYv4qlk8E[15:0], 1'b0}; assign r4JngA0ZVhEElGRZci9fohF = n0J4kP9YDHfDkhTNLn56dJ[15:0]; assign UpDw6anZs0bMPETxgXld9F = ({d8074IV5GByVrE9OuVeZYRF[16], d8074IV5GByVrE9OuVeZYRF[16:1]}) + $signed({1'b0, d8074IV5GByVrE9OuVeZYRF[0]}); assign b31KhkrKeVwOtEcPIkvs3 = UpDw6anZs0bMPETxgXld9F >>> 8'd1; assign Lcbc8UkQ7CVMIZTyIGqp7G = {b31KhkrKeVwOtEcPIkvs3[15:0], 1'b0}; assign a8xx20Fc5nKc8DbqSwNBuB = Lcbc8UkQ7CVMIZTyIGqp7G[15:0]; jtna8GP2YDGIaNOtv552aH KanolXBe3NA59HrsbrFCEG (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .pCWATI9lTIGbmXTtLuLAGB(pCWATI9lTIGbmXTtLuLAGB), .mgknRxAcgFrHqTt5CZvnSF(mgknRxAcgFrHqTt5CZvnSF), .sCFM4WicR6deeSAdSwumP(sCFM4WicR6deeSAdSwumP), .BKNY6GzA6oGZumjzTATycD(BKNY6GzA6oGZumjzTATycD), .uUcj3UAzjmPW47yNyzbT8C(uUcj3UAzjmPW47yNyzbT8C), .uwZv0qzQLi0MDBWLWzKuAG(uwZv0qzQLi0MDBWLWzKuAG), .n65LdbEr6NMNaEFcjX8Fh6F(n65LdbEr6NMNaEFcjX8Fh6F), .x9j7a5gok64zzNKnvdJNnE(x9j7a5gok64zzNKnvdJNnE), .bPL0FcLvoxhO0amTUOV9QC(bPL0FcLvoxhO0amTUOV9QC), .r4JngA0ZVhEElGRZci9fohF(r4JngA0ZVhEElGRZci9fohF), .a8xx20Fc5nKc8DbqSwNBuB(a8xx20Fc5nKc8DbqSwNBuB), .vLT6ef7BJliTDpt4k5jqF(vLT6ef7BJliTDpt4k5jqF), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .N2ZdE4zLlq5uRV4rcE2wdE(N2ZdE4zLlq5uRV4rcE2wdE), .iOhy3XYM3su7ndksftfCZG(iOhy3XYM3su7ndksftfCZG), .AECH0r3KnKo0RJFepDhYUD(AECH0r3KnKo0RJFepDhYUD), .twcuYIJzeZMBjyHmZ1FZDD(twcuYIJzeZMBjyHmZ1FZDD), .t30W3eeadZl9O9RnQCafyED(t30W3eeadZl9O9RnQCafyED), .flGpcmOyc38fKmqiV5eQvF(flGpcmOyc38fKmqiV5eQvF) ); endmodule