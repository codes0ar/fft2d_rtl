`timescale 1 ns / 1 ns module IWIdafyrOBWRPUGK17dNTF (v04pHKxyc2sPW047bbyUgE, JAMOfrNHxGSYDF0urqkLN, h4h0SDZC9CQgXKPbimISL3, b0pPxQrhAhYENzTiTGGny5G, jQKNLtXo0Dqi6Vn3Jy2niG, rosLsgtHKD6hJ64eM2pegF, j71O4t3Nm1w5MRqcbOUNtHF, DVmjaezJpTmh9E1RX58vDE, c50jzfprXP85SKSfjge64NC, s7ASYYS329kRVgP7KY37Y); input v04pHKxyc2sPW047bbyUgE; input JAMOfrNHxGSYDF0urqkLN; input [31:0] h4h0SDZC9CQgXKPbimISL3; input [31:0] b0pPxQrhAhYENzTiTGGny5G; input [31:0] jQKNLtXo0Dqi6Vn3Jy2niG; input [31:0] rosLsgtHKD6hJ64eM2pegF; output [15:0] j71O4t3Nm1w5MRqcbOUNtHF; output [15:0] DVmjaezJpTmh9E1RX58vDE; output [15:0] c50jzfprXP85SKSfjge64NC; output [15:0] s7ASYYS329kRVgP7KY37Y; wire [31:0] d2oEus6jJ0McV6ih95Y1AG; wire [1:0] Y8nU1xjYWVI5dgYrgIlsCE; wire igWwj37zoLbvMLlrefWxbF; wire PtqvgNqZpdLWxF206ad9XC; reg Td50TMNbpGWZYlXbqSVvTG; wire [1:0] f57E5i0241V1QEgB58U5YC; reg [1:0] htY8XTFJI2P1kmv6r9UdwG; wire [3:0] mAB2T9yHc4paNxEah9oqhC; wire [2:0] KhlHtRMHix8XvnicPL5XdC; wire [4:0] lFIFc1FMCEhdqlYwYW5oSD; wire [3:0] OP66o1rkZm1IVPqs42DN1C; reg [31:0] p9JdL74lJmHuomPqcevLHkB; wire [3:0] RraIPFfLtZsHXCwvliBhwH; wire X1dRLKXI3e3fN1rBDqxex; wire [1:0] WN8EiF2jALV8OH7W7KXXaG; reg [1:0] OAnPRhXN1f3PXR2YrHATCE; wire [3:0] bj4j66oAvfSpNoFLxGto1G; wire [3:0] jZJyU4ZP4ChZ5K7R8RriDE; reg [3:0] aIuu8srO6WIrizhN08OyGG; wire [5:0] la6NpbM3xhaAGZJpg3nLdG; wire [3:0] UAlS8hgEMaTiqrIEBR7P8D; wire [6:0] DB14wLF62mIfBaTI6vec6B; wire [5:0] Uf33riUqPe3QbDaMY9cxIE; reg [31:0] EVGDcYjDYMyphmfUWLd40D; wire [5:0] Ir5J1cq3X4AtmuV2rRCWJE; wire IfNgpXh3L8PgtuQ9riD96F; wire [2:0] rjTlAhUbkx4xhnY4CEQzSE; reg [2:0] Bb4Fv4CfcqYV9v1KrOFClE; wire [5:0] QBdSjsMcWKRY5gwAzbQLsH; wire [5:0] SxeI6Ebz4W3cAlBHX6N7HE; reg [5:0] a8prI6r0sJOb3uF5oZRDzvE; wire [7:0] f4gekvhdG5D2vtDRQuIsRWD; wire [4:0] HlCg528B0DhdId48qwIzID; wire [8:0] DdWFbmNZw3i61r2Flc3lJG; wire [7:0] C1ig1Tdqfa5ultBNsDcUCH; reg [31:0] RRY6uI32JPF7cgRt2ALKpD; wire [7:0] gMvZmbcqZ0DqgJ5sO7TczG; wire WPfmCIzxCRH3PoV577VFZ; wire [3:0] mIsPzyrzh6zMIEjXAztfSH; reg [3:0] W6W5MbHcLxMQiocqir3EcD; wire [7:0] b6B3OCDRqPO9Qa8fvVfkrL; wire [7:0] c0V0PWcNTcAtWfHHZo9oCB; reg [7:0] fCoWIZZx9VblaWmYgt13x; wire [9:0] btCYaoeB2JmWOR056EcY2C; wire [5:0] IgY2MGVmpmzbfdJvodzhYH; wire [10:0] x2qOSwxaMdgo7eci0FxvvcF; wire [9:0] baKrdskhfkPzPlkAHW54rF; reg [31:0] JnW70VzeuX4yEHMB8XIxSE; wire [9:0] p3SL7wYX8SBQnC0oYVuIuHF; wire q48UwMWOiN7vMKVlbAH62tG; wire [4:0] xTGR6ce6S4BzV4dkYyod4F; reg [4:0] jXOqwspdsCISwsGhcWqtUE; wire [9:0] fkhBlawaiECm3AKyJOvEc; wire [9:0] QDLMg0wJNF3uVvsVP11Se; reg [9:0] kfyELMjsnnzaUx6iYLK1a; wire [11:0] j3mLQ1yo2zmp8dnGzKOW5qB; wire [6:0] H5Q1sQZfYTS1fDeRqymzvG; wire [12:0] i7x1l0whvlbCztZ8yv9iwE; wire [11:0] ztLkXaVGX3w4pEn1xeRqMC; reg [31:0] rMhu2oApltCVSYS5itmY0C; wire [11:0] r46CEAiCE4Ch2WNWkeHtNeF; wire PloSd07HvtUIeQYlow2DsD; wire [5:0] wm9pXs3ggIACgFF4VQ65zG; reg [5:0] YfPairRXLNNVGttdcC4jHC; wire [11:0] actzjOg0aKNbyOOWNABa6F; wire [11:0] l0kGuUM557NseEtaykZ1TID; reg [11:0] wBLoEXjrUx0g620zErfyIH; wire [13:0] jARRiz24LDX5CAkjjvpbMC; wire [7:0] cOqqXZggK8lV63HuJIDU6C; wire [14:0] g03PW5Zn8wGm996TsM3OlSG; wire [13:0] seXC0DlX19Qu2W9b6laBkF; reg [31:0] YuoRtO5uahqj9k1hlroeUD; wire [13:0] VJtd7Fl5sWCBbwZ7zVkiAH; wire DFiuspHBeirfq1ZvvofTRC; wire [6:0] ym9Sp6nhcDPOiwj0UyGXsC; reg [6:0] zQQJr5Rr8Ek603tPKykxHC; wire [13:0] P1SxQfGkK55cR5k1YisfzE; wire [13:0] tp0Xxl65VoHaM4O6FDb2N; reg [13:0] toUJwGxo7JfW2EzqeaegqD; wire [15:0] hqJrTgFxozMyPx7LnmLBzE; wire [8:0] i3H4mRdiwOgMnPaGpxPykE; wire [16:0] IbH5QT2AXNs8KsoyD12ZfE; wire [15:0] V1kZ7bFxQFV1KrNlMFxWYG; reg [31:0] vAj4ixajCquQJTqGQyxOnB; wire [15:0] O219BqtpHO98GKSgKS8BpE; wire FTmP9v6IJWTPVZpRmGRtIF; wire [7:0] pv1WByjbGdV1OSiqH0ksnC; reg [7:0] DfmgsE3iMkzCsirhmlRDSH; wire [15:0] x40VeLX7J3a3tphEEkOgR2D; wire [15:0] n6crFALdZyJcOXZ3tAFGjWE; reg [15:0] q72w2glJ0iF1fL3kkboMy5C; wire [17:0] eUkkETd043d2fZQk8jDNbG; wire [9:0] ctWCGk8tDhNhqjRiNbiT8G; wire [18:0] jtIl02WJwApYjH6zHw0ps; wire [17:0] aEmD7oGZhl9CNV3Ln3b9jD; reg [31:0] u2ZdQtNDigVBNNBtq7C1PFC; wire [17:0] xUhkT9IaYCKujHljsYB4WB; wire aEXdj8byA7uSgyb9LhSHuH; wire [8:0] Yw6DjbSH20VSb4AH6J2ZW; reg [8:0] VlHUymZGBDkWniRKHnXeoE; wire [17:0] BmC7Waj3h156ApBRR8vBkB; wire [17:0] e6y0zTjYMJQBzfcOI5kwLeC; reg [17:0] goHRzycDTV9MFT2FCIUeIF; wire [19:0] QLgRzXPFcx5iBqm0rMhzn; wire [10:0] xbtGwTj2py2rKQx3DwaqsH; wire [20:0] l5Svt4GkcCOLXXQwBiRIcD; wire [19:0] wCUr9vYed0L827ZSFIusEB; reg [31:0] yI0NKYDzTZw44KqJ9a3zC; wire [19:0] bkWNTMVtSZYFA4nZXmoiEG; wire vlYCGljOoPPGkfFDbGHWcC; wire [9:0] SZm8Zt2WiFh8VGkrN5GsuC; reg [9:0] e56HDsGesAEqHwWeqzouMF; wire [19:0] zLl2QCAAjWMixlTOkaGHiE; wire [19:0] PcExrzPwT7phvvgF45pQHH; reg [19:0] Wz90RhDyGBtEdtGrJ0VTZF; wire [21:0] s2ByO9sLopwaaKB3OlviZB; wire [11:0] SRZlivglW4iODt3ZWa6YAB; wire [22:0] mTVvj9euDcz3QKkAdcmZOD; wire [21:0] ay59snlUFLNfqFr9K8OyMB; reg [31:0] VrDvujAzBpk1JUnt3i3jrD; wire [21:0] nXG6pKWoysTLlamoZb1kUC; wire FVZq6SQWJqDew38uj3ZwuF; wire [10:0] UJGgN0K4zoVMt8OzpDRhbB; reg [10:0] ElZOyt1VjSkVNH6qpuxaXG; wire [21:0] w0u8eyeEsFecynkh04cF1lC; wire [21:0] WXHkYoAaBaLUFbVOCc8VxD; reg [21:0] pNjnAf3CRLybq0T318tpZB; wire [23:0] pUZF40VeZ6xEJvpR7Es8FG; wire [12:0] CZy9D9fjHBHcfkgtp0KTFH; wire [24:0] kLW7ETLJg3f0fhJvPfzamC; wire [23:0] jV8kLyXAcS3FCyqURyzmO; reg [31:0] iLdfuowoyk1MtRrU15MG4C; wire [23:0] q9f5spD683cNlZnQf56m4ZE; wire qE7EncjwDfib2QclnYwSgG; wire [11:0] PPmIvwimSHZwNXz56Jo5FF; reg [11:0] s7H3AIDyv88anihczWgA1F; wire [23:0] fjwwR4v4yEuDBPgyT1rTBE; wire [23:0] JRbiQknn0l3SAzJguSaDIE; reg [23:0] ebaB1Kw2OvZfbCMRd7RH4G; wire [25:0] WOq3F3uShD744l8tfCN3PC; wire [13:0] te9YCAmyrsrdkIOdNQ10YB; wire [26:0] r0mlnEduB1ta4alefYkcSzF; wire [25:0] chc7OKgA3bugXJCo3yas7F; reg [31:0] lEZvI5hvOIId49rKN6EG9B; wire [25:0] d4IpN7AeFzlW8PIZDtHBNhH; wire kdK0vZeghYKX1pPI7TOLUG; wire [12:0] vIkIEBTGTAhgY525Xqzf1E; reg [12:0] Igu3qoayK7OqaCOGUvR5mH; wire [25:0] uR89cXy8xlRQIE7YbWSVVF; wire [25:0] jWK6QZgHeyt3ftPSKbIyaD; reg [25:0] I9gVg5rOTUbEKRzS4CERmD; wire [27:0] UTCgRY29pVn3brpE5SMH2C; wire [14:0] v43le787IqXWHekLEH8sc1F; wire [28:0] ERrwsqMxpQKfcAVllHsC; wire [27:0] NztI2AQnSAdBX3RAcWFzi; reg [31:0] nY5HJQdvwbdw1Z09MGQJdD; wire [27:0] ZH59np0e4GT0PI42ZDK96D; wire qvx4HYpxmuqVBKosKL9nDF; wire [13:0] vXQqwFz0Mq5pyOl5hUGpTE; reg [13:0] XSv77atgil9CALLij3LDU; wire [27:0] fqeYT46R9tLTDvWKi4sZDC; wire [27:0] FQVTrSjADBrb3DyvHSAwpC; reg [27:0] k2Wyo4gBkJTLcHbPeag55GC; wire [29:0] bb45jO7OrRC3XbD8zJ6puE; wire [15:0] XXiXbfRxJuy8atUhokFqtC; wire [30:0] UW4b3bm76Bs6tI3IYkPZIE; wire [29:0] q55ENw2wkQaVRklvIu1LrF; reg [31:0] aJrV9N3G9wp8U0g9mfcyX; wire [29:0] ZYrtxtrqxr2hmg5PKUYcOG; wire X1QJVAhYCy1C1RlcRQ7ehC; wire [14:0] cLzalZ4N3AQH17rH3HxvHG; reg [14:0] FoKnmJHxBvoWITgnEM5uGB; wire [29:0] u4MPAwPCLIAgQPn96oG4E2C; wire [29:0] muL6drwYusIoOSLLD6cQME; reg [29:0] ECSbb2HpHz8MkgOToIfkRB; wire [31:0] pUbtxeEGlqbH77tEidOseF; wire [16:0] OBIn9RfqwS76ifr6ctbJcC; wire [32:0] Vd09OCdvDhHzYbNi8eFYqD; wire [31:0] x9dWBNZVozdT9sZOUOShSwE; reg [31:0] c1Fi1DCmwETWogyXFP0luXH; wire BQlKwJMG1iIAM1sM8WOwZD; wire [15:0] U6NVSwrrDlIXWmZMGhGnGF; reg [15:0] CNCrh0XltTO38hUhsOK89E; reg [15:0] tuyMU89x2cRtnHZbS629ED [0:1]; wire [15:0] X4jT0JtvhLt1PtInljBofC [0:1]; wire [15:0] FTPlQQTDuHArhica0zG5YE; wire [15:0] ztGXs97JmxTgacz6ch5gZB; wire [31:0] kilI6xSQxSJzoqPMjerk6G; wire [1:0] FbKbMjw44CL9zGZx7WXzGF; wire fB6UnuVq9iLH8XGHOxxXZD; wire UPTJ0KHCAkQKe7namSEKjC; reg YWY1tbo2DIf9KVzn8BwzCG; wire [1:0] z1nwdQwUNbMUELLx9AUfwkH; reg [1:0] MEBenkOBGLeR7FTQrrn3MD; wire [3:0] O6EltwTicLhBoBnh9C7QlF; wire [2:0] WDqWbhmj05r4Wjj5vIY3CE; wire [4:0] cxg6xJXOtsYvHf3YKjaqmH; wire [3:0] vzZzLR6yNvm5R3q77DDCBG; reg [31:0] ecTpLKJNtox43CqRvB7TqH; wire [3:0] YX0TWRD0dHUDqZu2WRc64C; wire FCe1MyFX72qFVD3Hy9hPUE; wire [1:0] j6CDlg9BLVqvfP3aItxlu6G; reg [1:0] wEKIGBrNcPO2iCCXrGUIu; wire [3:0] d3qzATGoyxtZcYJcgfDfbeH; wire [3:0] nOloqK6lS4ZdzwyM1eUzUB; reg [3:0] wpq9P4PBi8CGLKpUN7fWZB; wire [5:0] o65FJTz0B7IXjYcgfpVqSZB; wire [3:0] C47tZ0C1xf5jlTyv6MLJdF; wire [6:0] lzW16GgG5bSiyHby6MJi7F; wire [5:0] o8P0gThAuIs85SmAegMaBdC; reg [31:0] NKytYt7HRGpr10Je7y72bD; wire [5:0] r5YWTZbOV1ZMPt3R1VWQsEF; wire claoCCs3pNDgkEZUVS4BEC; wire [2:0] QKjfaK9XJfQuzgSPqcdG; reg [2:0] PVfspm0nrz7RTrj71zZK2E; wire [5:0] bcdChZWFB9riH389qHJhvE; wire [5:0] JT69Ak8v7evsLSjX2WQmM; reg [5:0] t9R7A1peR6CuzTzZAm3HwC; wire [7:0] QOFovA9T9qIZcEqTAPhtOF; wire [4:0] iar9KCTPqGuEmE9kiyh5vE; wire [8:0] gCZzU6M0PYvvj8GKTwHOiG; wire [7:0] f1zvQhGH1CAcbvWG7t74yHC; reg [31:0] Z4I0KdM2JVi87xjTMS96pG; wire [7:0] nvyG06fFyy1jvHC47zz9RB; wire cHWq2LRdov1nvfvvjvk3TG; wire [3:0] l1XFmcvlNKvaQmQZV9JV9jF; reg [3:0] EokQF3Q771FYsuXM046eTE; wire [7:0] DFG5jHCJODhySug0Ml3hXC; wire [7:0] nqmUVeMYCM820YVZt5ilzG; reg [7:0] f0Pv94BMpwnCMzWcufXc6hF; wire [9:0] KbzFknNUACxVWcnzlxJfPH; wire [5:0] vQdMrvqDo8qF2kLKQ7AeXC; wire [10:0] MmjkPa4HYQ1KxOVnGr5TS; wire [9:0] KiJFVa7Kln3PVycUSEnQNG; reg [31:0] npDxBmN6dOapdh7YCQNR6E; wire [9:0] l9uTQkxnOKF0VsYALlWDi; wire df9yw7V8ETyRFsW0D9NBP; wire [4:0] x1EQwZFojLp1LYxIXBaNWE; reg [4:0] upGPDbRFmGJ0jGUoSFSlo; wire [9:0] scXDy9YYbNjMkzYu9H6NVC; wire [9:0] uZFlhddYpWdV2PRdQqigiG; reg [9:0] SYr8j8M72olItx5mxZg3Y; wire [11:0] ciJx9JM6wpMOOlrHHiFDNF; wire [6:0] S2BiHHBn9DfCYxiINFX69C; wire [12:0] A5VMUTy53cH6e5xVrTmqs; wire [11:0] dp2CW66DVlddH12FzsbYtB; reg [31:0] LXl9oQE5X1sFOi0vAmIARG; wire [11:0] TaL4eG7ansmqPnA9GOrj7B; wire ovy3LStQ9NhYK0h8Fs3GuF; wire [5:0] nFECnxinHyxo8igKFGptnB; reg [5:0] QVb00VBEtaVfpEONJrgsrD; wire [11:0] i8Q2fmoBrZj5QeOKDTy7OXC; wire [11:0] aCdbqb3Z1RZUA24wJhmb8D; reg [11:0] d8keq4sOv6FPsVBE0yF3SNH; wire [13:0] u5OcuPukOTULEzZHTQa5jE; wire [7:0] pnxSnkOhYHGvcrejMZZzGD; wire [14:0] pc28A478dggU3B9LCjrwKH; wire [13:0] Gx4uCMMDMcZkPFg5X7j67C; reg [31:0] VyfaXsLYCMGgAglyPOPl1C; wire [13:0] Z2TjolWsiqSfSlQUx9priB; wire vHqd7R6RAG8NCgLXFiRG5C; wire [6:0] j2LzkDa3ilhqsCEzuuaMJF; reg [6:0] d8vwhmLzwzph5ZWCJmi6ErG; wire [13:0] POoNYqus4WpIeJLkV05T5D; wire [13:0] Rz1A4aD1tARfsL4hWRkGuC; reg [13:0] zE0XGJgmBnFBVyzADLIUtH; wire [15:0] f7vtVkzvkHLoKRQDBqXTbID; wire [8:0] xtUeqmfA0OlZnZC5um4zvE; wire [16:0] l1Zuzf5TzQSJzUw3Msm6HJB; wire [15:0] COlOv7R0Bf2iQD98SJNBZG; reg [31:0] P6kiEiTnuWYRUMrtGnBCNE; wire [15:0] xbOF64W9Ar4Lqlq1uimKrD; wire j7fDTHKDIw1b9ho08HQpp7E; wire [7:0] as3iWC3h2hgaDUNBaZqgv; reg [7:0] UjnjfhzZkOwIVGTyKJXtgB; wire [15:0] p5quEV42RCn3OtXuG3mHSvH; wire [15:0] kbuD4rfjFj3gUIhRcx2cdG; reg [15:0] QejN3kgI3Jo6juzY8hBlyE; wire [17:0] IeHprHWybCEsl7WYUcFGsD; wire [9:0] JIAufNDlaR5FZG2gmjhTkC; wire [18:0] ru0nteK8qxRvyWKiCzOgyF; wire [17:0] o4ibQVfuhBHTF5NDhAQ1fKD; reg [31:0] RtvTaElUgdpBmXzJb0yJKD; wire [17:0] MyltTFSsXFeoPojqyAjON; wire hXEYb4xQxcywPjqLBUEGgD; wire [8:0] p41v0Mk0HADN0WDJBhiMxfC; reg [8:0] ffsa6OEyoM0DX4OPlTzw8C; wire [17:0] nj7Uorw3TSz9rKxp2igQEC; wire [17:0] kmD6Ilrh464BCBLVMn4VbE; reg [17:0] kfbQPocRbakJ21Bwqsv0i; wire [19:0] Iab7HeJSQoSgUz7RuhVazF; wire [10:0] jJ5plnxESkvDaAL3rZt2LB; wire [20:0] QEYaVcLKCNUVOqER9xXxWC; wire [19:0] pt5fnF9KyMic6eq7rU7gqD; reg [31:0] hrT2I9W8UAX8lkCh9HwCyC; wire [19:0] cfe4isuXwwohZOaspwNnNG; wire xJZJ529nCjQslckQHtmxZH; wire [9:0] j7nAYb6dlFCqOFMxfcVd7QH; reg [9:0] JHUut6Rpogqw8E9skISIeG; wire [19:0] TE4W5J0afB9JODLAQ10TQF; wire [19:0] e8QGmucX9ku7ugMNMP8ZiS; reg [19:0] gpMM7ieMx4QRfhCV7UZauE; wire [21:0] OUglDJO4thns7zNL28NuxG; wire [11:0] C7tDtgXgfSxjvHdfE2p2hD; wire [22:0] CyNDnUuxJcv2BmXf9rWncE; wire [21:0] MEVPG7Vi3Dy7JBBjWyUNc; reg [31:0] azzFEVo2AvUNoNmYWBwoqH; wire [21:0] eeRMcqFduj2oNy3g1HVxSC; wire jz1BZADe0coZodBEtJnz4C; wire [10:0] IwuuD2S9yNrHHdvvAG5YUH; reg [10:0] imCuL1FFwqq4jnPaCveL8E; wire [21:0] k2ck0YJnFDXHpMedhgr9qRD; wire [21:0] sDVB7xEtvbOFj8Ui2bnoQE; reg [21:0] JVzqyten1mMc4Z5uvlfZDE; wire [23:0] b88drpPnD2VtwJtiEYRFQsF; wire [12:0] qKdAaZR9hfVY5g9WEB9evF; wire [24:0] bswyonmpcfI0PoIt3aDSnF; wire [23:0] BzfSkcRvRiID6B853Sk1fE; reg [31:0] m2hoy362oakremk4ykeoJB; wire [23:0] a2E5bq4xG9P8XECnOWVSMB; wire s3Q2hbnFvcjqlvgMHyoBJE; wire [11:0] bZEiDJSctoVjsoXa259StH; reg [11:0] eDBMOFTBb83n7sEEEKLXq; wire [23:0] hvkiJvP1syVDuE7eNoNFYF; wire [23:0] cm0e9uh59eoFN2OUKptdvC; reg [23:0] EtkP3DOGdC8t6olD8mZndB; wire [25:0] iWvOu13ViXR7sawgPT1FjC; wire [13:0] FCMxV8HogSFueL98F2gNZB; wire [26:0] OqbQk3ID7Nz1GCGU2AjVl; wire [25:0] mCdg923NHIP5asuuf0W2lH; reg [31:0] UWcy8pW199vG0VtRCBW2KG; wire [25:0] ioSpbvR6GmIfKRjNpsh2bF; wire WX4RpTNKBdQSVBqSWlRVFH; wire [12:0] T49urcBbEEYXRINyVdZulH; reg [12:0] e1HEl1XlshKTotIEunk6hl; wire [25:0] w7VJdxjubq01SlsqGHlxfG; wire [25:0] tTlljYwJT4O5u3alzMe2wE; reg [25:0] QPW8GtDQnJ7lqvnVJpijxF; wire [27:0] X8nA6uSQZbaymM4A1xITNC; wire [14:0] iRy6kU8Izv9CM66zbzdb5E; wire [28:0] KP1LyZ1AFIuavnuOnBw1VF; wire [27:0] M6VKmyjZQOZXGkAKz1YjmE; reg [31:0] Aj7pH4hZbnjAUjVZDj9vFB; wire [27:0] DwBwYHrLgg9kBDz3J9ELdB; wire v4mEf9URPRBLqIECbXnBDH; wire [13:0] NKWf6OMVvpkOpk9VSSgyRD; reg [13:0] pQouavJJCwsKCEciQhrK3E; wire [27:0] bEAowsULkF3zy5hFKpiuSG; wire [27:0] yJA4o0iAYXBOPsUCeScNfC; reg [27:0] IeN8KMSMvMg9IHSLo9n8DD; wire [29:0] zJ4HWiLEv2XMiMoWf7FLPF; wire [15:0] AVFpT7Ib2pO9YuXeN5BZ7G; wire [30:0] f7EfvG50GJ7jqsywvc9ALC; wire [29:0] i0wZxrICRhlPz2FiwtdU8D; reg [31:0] Teq2Ch748yHVvAT4uGB2FG; wire [29:0] u5WmpPBQNytMuE3KlJIOpi; wire o3K5Quha1VLfPYfrjqgd2GC; wire [14:0] i7el1SwQPx2WBbyDGEvo0HE; reg [14:0] KOx599mHUoBor0KqJHxFwD; wire [29:0] faBh6P2w0PfMFOrrdKqngC; wire [29:0] Hh9HmtirCWU1zK1p4lc56F; reg [29:0] BqdWvf3iIjFaDgt9oYSkhG; wire [31:0] SfhLiBMyxkjp1mCnRxW8FF; wire [16:0] BsKpUAswevf1juloThWu8D; wire [32:0] RSGrktqBvyzhNztToycF6C; wire [31:0] a3rKmat8RqcNJsLf5q2n3lF; reg [31:0] rIrurMdcINDtP7R4SI48FC; wire TIXiaddILO7mGZ5fWGjDCG; wire [15:0] q65RX0Z30mhM7iJaeWaDrB; reg [15:0] huOSY5XC1YM0brxFNzDqbH; reg [15:0] a0r0hzxzkyJf9emryhMzNH [0:1]; wire [15:0] mSur73tREBGM65xgjFu23D [0:1]; wire [15:0] FbFmmmgZQfWceRTyvEh1XD; wire [15:0] rli8whUrHAa4gMtjCDSb8G; wire [31:0] D3zFB0T3BdpEDXphszsGdB; wire [1:0] CbG6VEOygHZYUZzB34fCPD; wire LRYct7GPXlUHbsVioc1vsC; wire O5ZhenpM9MNYjlC37pcmaB; reg VFANHQZIGPAY7b4qkN3UmC; wire [1:0] wPuizGWKwJU15dBqzdZrBD; reg [1:0] mqahydaC3BSODO8RxqH5PB; wire [3:0] VBO1aVfkto7xu4QNiqWIZE; wire [2:0] LdC0oEIcEn2u37BATOVquC; wire [4:0] kI3sx5pDEv3shi2CwtDowE; wire [3:0] PHhhAthYaDH0mmviJi8guB; reg [31:0] aT9efCDUWqkTFzkLh62zcE; wire [3:0] UNAFAbTORoRqY4QDbHcJqG; wire AdwV6s2RyWCMBpwC2HwLhF; wire [1:0] aBGGSCfHl2skiiW7NMSRqH; reg [1:0] UIRrrD9huSjdHRzMx7sndE; wire [3:0] ws9KmMi5xRwv9SWSpHlEjG; wire [3:0] BhAtwwns2SYFGkylFXi8BB; reg [3:0] bFIpPSFT8qi1DFuaWqyHtF; wire [5:0] V5pkjBsnPThxfTE1IZqGDB; wire [3:0] GgVTSIzPhN9ZDNsuxXlotF; wire [6:0] sPR4NMAZgx7B4yl8mD6wTF; wire [5:0] NRJsb1CWMjRlknrudNj0vC; reg [31:0] d1GIPVaPfFgcgiwAjKvy8SG; wire [5:0] jjj0aH2qdZsn98a0jCTomE; wire rv3m1T8mIpqw1vC5V1KXZD; wire [2:0] IiAS0qAOkfTGhzWxyd94bB; reg [2:0] NR1xVi9KX174l32cXe7IJE; wire [5:0] lm4lGUUMg60sZsVKf4JVgB; wire [5:0] ivLtaKVVFqPbuQPRlcJpyD; reg [5:0] n7foXfKUGohH9shaofl43E; wire [7:0] BS57yRSQtZPyqi5Bnq9psB; wire [4:0] bJL4EEMedVetHndvDEZV5B; wire [8:0] h1eiDNa2zA9F1HKjhzXOf8F; wire [7:0] N23SExOhay0JnnZmBL4yeF; reg [31:0] cVgZOzpOdguVRHYqjIhuk; wire [7:0] UeTfFS2ghyunTw4P5wojCH; wire r2aRRQzAghfWk6CnLQvNaED; wire [3:0] z0UZNzqu8Mq6paQqQqHK4UF; reg [3:0] XXo1SDyBQiak88sFppTsjF; wire [7:0] GY9QWHEBZRjto6a1NRA3iH; wire [7:0] zqHHk5KgIKVa1DwUKAqBXH; reg [7:0] n6lFBOQkulfdWipZ1B3mg; wire [9:0] LfqJxMx8aPdx9Tg8ZpQLDE; wire [5:0] ksNnbnFsGUzsj0zxQU3sKE; wire [10:0] a1iqvsOthb0rcqC3PKWRQDF; wire [9:0] YDcXhhOhmGwMKoHYiwexTC; reg [31:0] HA7EYu1tK22O9i8DfpQe9E; wire [9:0] kJiADoCkwzhBqxbx6PgBqG; wire NxDv9cBGuOcye1qdzN2ZbE; wire [4:0] fkCZV6cvbAqBisxRxI0dSE; reg [4:0] e0vzZybk8EaC0sU9yzfVEbH; wire [9:0] KX8K4bcTmgK9iJZ4tFToED; wire [9:0] kaGb2Rgb5TMNxVjGWXMVbC; reg [9:0] c5L411ATxQWGbO5OX1TqZgH; wire [11:0] iR44CzvnLIWQDJIT2Bh92; wire [6:0] ggosYHNjNRgTTSM9nJcDSD; wire [12:0] z8NqtohpOQLMO57InnmOb; wire [11:0] q31ojLkv58ZnYslUMTLzsC; reg [31:0] smVaYT3RjC4ThcTM7llQyF; wire [11:0] p4997dIwDfgVVzHbKtpv7QF; wire qZOy2qjQqYVt7j2rqbDCTG; wire [5:0] QoD3LztlGG71FSISslVviC; reg [5:0] phuPRYTWQCA8RK13saxVWH; wire [11:0] bZbQIJNhmFe85PbMpnosoE; wire [11:0] qtXfts89aIY4wmBLUXPOB; reg [11:0] NuscntgAE20ZaRiAV7hqxC; wire [13:0] kPLHo9hogSxDdfOl2CHNl; wire [7:0] t8xCnJCyFWgQ4D81QGbaPYD; wire [14:0] pQltLIbYG2q4aRwtQURJEH; wire [13:0] Lo0IPZ8YOZYiEHpLO42t; reg [31:0] x8T6JyOFCXgf5J8GjRm7OkG; wire [13:0] e9iuXqe8OquZNIsYKIaMIz; wire HDdk8UacCG1vTeipSM5kCG; wire [6:0] B6E15sMkwvf69CPgeXdeMD; reg [6:0] WgndoVXG1lvIDs49UGDJ6E; wire [13:0] pyOvyPa77c8LmSRqhL1NzC; wire [13:0] Pumm6kexkeR2FSC6LmP9s; reg [13:0] OVKm7tgpOSGLpjnZC3LTHE; wire [15:0] aU8NJptrwQ0dPQIyaGkVrF; wire [8:0] Js298tNl0lY511TfteNPUH; wire [16:0] fQjzw0fgAbUvXvStCKuH4F; wire [15:0] p8Ah8TzME5owYP5XfqJRi5C; reg [31:0] w9wFocuxSkWDmPJPkThqR; wire [15:0] SIrY8D5zdov6veAntRlukE; wire DDupKb1BKahfvyZFNYIkJG; wire [7:0] pmpGHYek38BzarQ3qCmQrH; reg [7:0] JNYY5yF3xZ1TK4lLNrmXEG; wire [15:0] v7Sqzflwbh5pKJBPCHTKDEG; wire [15:0] IDrfZ6G75w0b2Ygh3LfQqH; reg [15:0] Jddhqf0gqhZPY3wPFOoq0B; wire [17:0] n8scxI2E0ECdA36CQrpIbcF; wire [9:0] d7Y8ztVAPOhsm7hvfGhOi8B; wire [18:0] IowNApmWP2sledCgFHJxK; wire [17:0] Sg8Rlnypyf03avWXdcL1OG; reg [31:0] XIKIDtpbTSIlhPajFWHSwG; wire [17:0] pvJes4iUAsoX3Tn6rjCtoB; wire u9XFbiauz7fSkqkXqpsNWG; wire [8:0] w2kjxMWJYgH9lTQZFzFa1; reg [8:0] a2rtoOfWEDzPhJ99mgT6QC; wire [17:0] wWFbZBQIqqnL6q7blY0Yb; wire [17:0] QIgCUQ7mCaVPNoxTkCAy2B; reg [17:0] bZ0TC5wIi5iy30a4rNIkDH; wire [19:0] lBNV6ky8aHM84IPsYJR5n; wire [10:0] CncqyghSqUQTM1BqMCiVQD; wire [20:0] Jz4Rz7lGPIBJhH3PnjgUm; wire [19:0] AZ2r2El21cWt3ILZ6XvcTH; reg [31:0] rsQbmn4FST8xbRglSdx2gB; wire [19:0] iDasY7iIgz0v06oml0mB; wire n2bWPIO8uW8vas2OgVHEQG; wire [9:0] R6Vz9nbYsbvk5sgLGoA9gH; reg [9:0] wgs5gJPwk0LvUXsr88hTAE; wire [19:0] f8MC4kvmiJjXr0IW8cxs2JB; wire [19:0] gI1jgIcglDsIX7jWy9Max; reg [19:0] qg1fRXQtNbgVxdF6yoyREF; wire [21:0] T19dIaBYdTa9PZtZdWgMkD; wire [11:0] GP7CX1dPzFlgdxhmIe77IC; wire [22:0] ukHuAnhlCk8KBBDJvvXX5E; wire [21:0] WG8gzdLTcqsl8GywHjG9d; reg [31:0] n0NkQdqqnvMhDs423VLBKB; wire [21:0] sTeAyrqG3sAnFH0TEwCgCC; wire VFMMCmH313z9JCR3kquowE; wire [10:0] z9QhOFznxLqChUzhI5cK0jG; reg [10:0] DrSlN87zei4SgG4DNVrvDC; wire [21:0] f7JMRjTBsPaAUm0MdIgRtnD; wire [21:0] Xi3P8xPk5lz5vI0tMPsr6B; reg [21:0] f6nkTVOkasMPYCVdQ1t3RWB; wire [23:0] zjOnmfxOzwLbAed0PkfB2F; wire [12:0] IfZ4i8sgfnUgsLonllpv8B; wire [24:0] E5qxoP9J21gq2LElkgURED; wire [23:0] vAlvu2utX7HZnziQ9vOxcG; reg [31:0] m4y1ic6jtAcK6wabyszk2XG; wire [23:0] IcVjQXg4SRLKRiJxxXqZ8E; wire deQ1vqISll3LmEKYH0A7SB; wire [11:0] c7yDah4XfUadElmPskVmLyB; reg [11:0] Nw9XhYz9rDGSiYWFthwTjE; wire [23:0] JudNijS8FpWpflBOEYDLHG; wire [23:0] b5qQKAR0z8iaZSmFCHxUOB; reg [23:0] jTESx94Dd1T02ZzWeEVYcF; wire [25:0] MMf02FL20h69sCnNPkyTnG; wire [13:0] yBpiynqDUQkwe3RYNavApF; wire [26:0] NOUvhKrq6oFXDc4VWYTVdC; wire [25:0] gMtX3xfic7tHemznuopkOB; reg [31:0] j4Arti1lMtcMN8FLTYwnLD; wire [25:0] U2Fo3lJvtLBHW9ogfdvMME; wire hTRZGt3YI59beY9UH4p1hC; wire [12:0] jCWS9kN2uVkHBlJLgsj6kG; reg [12:0] j02zF9SZU2kTOSADrFEpciF; wire [25:0] c2ODxgHWlHLoVp7DmYQghEC; wire [25:0] VZAGPjw1JyEheBnEY0qxmH; reg [25:0] FEy2g40kN3tEW69WdAEGuB; wire [27:0] f7yOZ4lKvM8fXmfyUsACQD; wire [14:0] vgJ3Cr2LvuSOqY4k6A7uGE; wire [28:0] cUxMq6Y4mcjJgTtYxIGyAB; wire [27:0] xl28WnwOjU80W5ASAhe6dE; reg [31:0] KHqMKdR2LLNMgtSzPORlmC; wire [27:0] NUD6Q6W2pS2fgKUnNEVCgD; wire lg3UhZcdY7ALcP5blnn8XD; wire [13:0] zVMIcJdSJmTolQAvSVleTE; reg [13:0] kBBAFkyIMdTw9pxAjJ1PQE; wire [27:0] d7eCmZlCMqvmGdTJawNyWjG; wire [27:0] rIdmAf73ZEwrWcZ44F3tgH; reg [27:0] bpSKi6hivc4nH6E2zzIO0F; wire [29:0] jh5AUrSuZO8wqZbeaVRW2; wire [15:0] yhPwQJOLmQPtFG08fBKjl; wire [30:0] cyg0eXE4VhRBBjgceai4dC; wire [29:0] e29MWCdfscO1uEFKXjG5E; reg [31:0] I0k15e4Mqbps3RkfuTGQjB; wire [29:0] TMGATS9eD79sBvLQD4W6iG; wire WiFgj83PIvYCFc2yBQbeW; wire [14:0] a5WzJ7XQv96wNGYwcc9tqG; reg [14:0] ipdO2sWhLe9H5WGpausKI; wire [29:0] cIi6w7oMwXcWCEETgy8lPB; wire [29:0] JrtSMcosjxt3HtURicDP1D; reg [29:0] mEmXvk5JjuKgxmWiD2PTKB; wire [31:0] axcp60hEFY4m3CLm2qD0RF; wire [16:0] jkQbtWVNPA74tjUiciPhpD; wire [32:0] tLOPvPysS9xFrLzWomBlzG; wire [31:0] v4pxjsLZ10u8ylsW5IyGeD; reg [31:0] AU8kfu9Bk1j6iNF7JHgrNC; wire adhdaT5bCy3ZoSykpu78oH; wire [15:0] kmeXG1ZdV7nLMdzktaC88C; reg [15:0] oBIxcPTGR95iZNFbr4227G; reg [15:0] s16lp7vAtcFZ2wwPaIkgzB [0:1]; wire [15:0] QH69kVWWgj2WJadmvpUaPF [0:1]; wire [15:0] FS8ak02sQNsotNaSejJzOF; wire [15:0] s7iMbfZ00UZszqLEi06wYE; wire [31:0] YAPbE5XIglo6YQglskaaWD; wire [1:0] b4c80DCXt5syU5YZsPFg8fG; wire aeA4SROkYBwZ6Vg6wePll; wire VLU8KlCAVdk3z1akf8lgXG; reg b00qa2rJFIB1ZMqONGFopXG; wire [1:0] xmRFmcImcIZ7hAGSB5Bu8E; reg [1:0] SKbN7GhZfEspFZRKIkIVmF; wire [3:0] Js5jS7mG04lv6SG081bBdD; wire [2:0] n1zMPjaeIWPwBCg7gfpFRw; wire [4:0] JSVnqT7wQsMpSEZncqnKU; wire [3:0] d8YQiHX7vIPrjtzcNsFfqUC; reg [31:0] PkXpzwBbQLQYvzhTqlk7wB; wire [3:0] w7Sh4wi1uZ8tdPQjGm2IyBB; wire JIk51ZYgI4bjmkaz1s3ocD; wire [1:0] p5vFo8g1m0abgHiHdIbMIB; reg [1:0] nNsb6XV1QdVOT8po6E0QRC; wire [3:0] f2eRR8CFkJiACbGc7JLrHC; wire [3:0] m2es1PMsJ2xQuYLiPnHr1; reg [3:0] UGlnA3qCFkn9R10JNKEmWB; wire [5:0] f7i6sgURXoacv9zlCx7k8pE; wire [3:0] gFnPRfLYr5mEttAuZT5TNG; wire [6:0] AFbX6YpTqq1eBEyQFqseMC; wire [5:0] qqZdHvncdEpi1f3UX3FiLH; reg [31:0] Pz7nVzONTu3jrA61HPdb5G; wire [5:0] cr5TMAj7bawp4OzGhelvYC; wire uSBJDL0TF4CJ5LqsokDLtC; wire [2:0] FDrOrbrGZpLR2snFBNYfgG; reg [2:0] y1AuRFIyn548BXgwQF0sZdE; wire [5:0] U6ZX5GALoV26phzqBZLxwB; wire [5:0] lEpIUGd5Cr0vd5frOPY3ZB; reg [5:0] Y1kJ6m5YlbS5HZjCnkaC1D; wire [7:0] OsCJQX96BJolsZ5d0oBzoG; wire [4:0] MXb346opbIN11K8xrTYv0F; wire [8:0] JiuDBTKkk3DmNTKhQeVyEE; wire [7:0] cepH0TZ1Fi8TpQGwHx2WYE; reg [31:0] cUOLCqZop1yocpR9PH5jiF; wire [7:0] Y8QYTUsOLW2ORrnUf75Vg; wire mRBRsCt0Pgu3ZY8PRCi0oD; wire [3:0] n4tG0JS2MvMz1aVTykyRDpD; reg [3:0] CI6B2HVMFRzDx37oEWjIuE; wire [7:0] VSMVYe1a2T37zL1SHKrC2G; wire [7:0] w2M0mYanih9pVwcHbeGmhkC; reg [7:0] x08SSTqzuST0npo22yvHD1; wire [9:0] NrGTCqt9rkin8JxxJzivMC; wire [5:0] sMUm3XDWkY9euUemzzSHsD; wire [10:0] qjrpTJyWev1g925QNDAW1F; wire [9:0] SFmRqM1SKlq0XxdjenL8yC; reg [31:0] darCJM0vPSpQ6IgQNZHgPC; wire [9:0] YQ3g2H8nF3dqmEyVDvXGRD; wire PSPwNHQ13FhdLM6OMJRHmB; wire [4:0] NQ4pAf9vZ8Xx4lGiiOXU6D; reg [4:0] sJ6GWhkNdag4yzDVnIXRZE; wire [9:0] ObGqdHNTbg4VcYpEbgQjKB; wire [9:0] DRHq6AFeMUbFXJu9ozWhfD; reg [9:0] aAlJVECF2UJ0il926uH1xF; wire [11:0] y1txMzBbEmvxmMKJpM7J1iB; wire [6:0] wSKM2kCYmT1b8JpcHR77rE; wire [12:0] p3FlB7G5wQcEKEanZhV9aF; wire [11:0] v4aA671Zjc8PT2J1KV8nzkD; reg [31:0] URZZIGLG4aIgBvyK6bwvuF; wire [11:0] q92Pz7xfru0n25cOdhefGB; wire nqCCuMllPTQCxAwb4BAHtF; wire [5:0] m2Xf3fQbkf2EKah6ia1rhrB; reg [5:0] DP1rxfHwjNcmCS5dP7UEvH; wire [11:0] In2u3aBla1oHkNHMApLKsH; wire [11:0] RhvWLtfm9kbIPah6Xmhz5B; reg [11:0] ulxawSs2t7mfLDUIwzjgMH; wire [13:0] QogFm8TTkYvdd1pOETS8GE; wire [7:0] odys5fwKXDkTPl2xGW5md; wire [14:0] jUoV3u5hOQ3V3P9X4L422G; wire [13:0] lKy8gFEyss6k09Lab0TIyD; reg [31:0] o9IXOBjy3eJadOxzwMZYCD; wire [13:0] afhwDwKsffj7ws30MIdif; wire gzAMKqGsdPMTGqF8e9aodB; wire [6:0] vMT5nzjGBRaywF0w7bpHnH; reg [6:0] kQOxLlINqlKIXn0R43wTvH; wire [13:0] GIyfilklKRkkteItBi4jVG; wire [13:0] cDG7Ga2x2ulXJ9HZ0kU6XE; reg [13:0] cOQeVrl2Kc2AaEV3A3SKVB; wire [15:0] oUr9Z0wSJ8NEbpWbUr40O; wire [8:0] v99YLq8JtK6czSdvv7sUwZH; wire [16:0] OlUTROE94KsCPuYIZdRVnD; wire [15:0] q2d5CtZFCBdgowZqGzc7c; reg [31:0] XMliVuWBVwOcOPEdVe2sbD; wire [15:0] H7HCojLu6xl0FDsspFgeF; wire V5HChjE9NVsTIubsNiixTD; wire [7:0] r0fdrd8QpMOua7OUDgRkvlE; reg [7:0] ziHkTpSLxytlkstnKqPgtD; wire [15:0] TrSsPsucRJCHZyiwqiAxYG; wire [15:0] Bbz9EGUOWN194RSqeY9vzE; reg [15:0] P41QmEa2IVlG6Gw1uNCuYC; wire [17:0] liAyj9i3OaG5qj3ww4zBjB; wire [9:0] yCyP1ziVlDiJpYzdd6YPVG; wire [18:0] arTIxO8ttVfgZOyW4PzlzC; wire [17:0] dCaoI2qtg6pmjm3MVxzJKH; reg [31:0] dCOpIGH8phIdHUSJlDSfvG; wire [17:0] oflUhi5A8v1YWG7yE5g8i; wire g93FJ0IBN4c66etyHmEs3zG; wire [8:0] OeVgNvqOmoHvuonJYQ60DE; reg [8:0] zQDpOsty76yxOjWPsK2jX; wire [17:0] OnMuHOtaSmv6vr0BtqpDUB; wire [17:0] h3EKSUN8gsftz7jQO1rdxBE; reg [17:0] Dgv0nOPwuFJGc4GAqTimbH; wire [19:0] woO6WUPEUZHhCxslCmpXsD; wire [10:0] n6flnvH1JRdcq5tHRAY4lC; wire [20:0] Y4ORnDxB7EutyM3R3AYoLF; wire [19:0] kpoCQdFe8llOB4VroSkRWB; reg [31:0] WpoaYGV1NzHQJMT5jm5HyC; wire [19:0] p5ZR7b2BqOcgrhqd260UTF; wire G44bIdnYp2VbJFdrHB9ZC; wire [9:0] ZWAF6ra3GkzT56Oefe3NLF; reg [9:0] ATgyH1zIQ4sJ6Hz7GqMsCF; wire [19:0] lIdXhiWJIC9ldEsDa0NXZE; wire [19:0] P90P58Xa7n44tjlKivSZ8; reg [19:0] gyufbtlPcbpsc3XTEswKdB; wire [21:0] H7hJJQFtPQpIus6wdn7lu; wire [11:0] jCUl3tPIcmmqDiSckg2hhD; wire [22:0] wIaIyn7lrKf0kblWE9XkjC; wire [21:0] fFumSIcnLnWln2qYLinPuE; reg [31:0] nRdqcvDbm319JQcsXwul4F; wire [21:0] m7vHNxrFnoDjp1IrlzZ9fQB; wire QYXTpn7JNO59MwFJCQmpxG; wire [10:0] Dx1qecvaNRk0C8Sp1BRC7E; reg [10:0] YJM4uTYV0GNEIq6Ts1WqdG; wire [21:0] u8NrYi3OMqbhK9yByGZs9PB; wire [21:0] rwO0PhKT8dAkniV0s365fH; reg [21:0] QEFCsmo4y0LLYuDoykR98B; wire [23:0] RX0sHsM1Nzw8rn3ouqfTE; wire [12:0] uiKvXhWqzaIyVELDYBl2pC; wire [24:0] VpP6fnKzcKN32HJtlCGIuD; wire [23:0] e3PfhueHdzlIuEVJBllUSi; reg [31:0] PQtoGuipN4OobbDKTpW4zB; wire [23:0] kvSoFz62JUu4jx44u4ZCsC; wire vg0CbYzueQThdby6EnMwrC; wire [11:0] gCzr56bCiioiPJ7vxpKGRE; reg [11:0] g1i4ElfCXQ9sMqQ8agpYlLC; wire [23:0] TrlkOR4z072dMOyjD8yJtE; wire [23:0] pDEdPRJUIcsUQQ8UmXGdJH; reg [23:0] s85203G8LCtqp2Q4Hln8eDD; wire [25:0] voKrZH4np5NWTctmsz4oFH; wire [13:0] e1Rl7kcQNObhKfOXtWutrG; wire [26:0] Taj7HNFKppS43yrU3qKE1B; wire [25:0] L3nPxZVh5u3VVA1rdbb4QC; reg [31:0] DqFCXgxzTWTDDQbslRF6E; wire [25:0] d3KDtpVH3H0bcfiybpzeSnB; wire sGiOEpItJbE2kz8n13WEwF; wire [12:0] zFwPpMKHPaoWNlMcn3Ooz; reg [12:0] L8G5zN2h3nNrCok5TCsJbE; wire [25:0] BOaYPwGg4vIF3dmZHl7rWE; wire [25:0] IJwTxkeWtn7iKzAUHVUPeH; reg [25:0] DXqu7TpZsKBJkGAUCIfEdB; wire [27:0] wxD3MMuIUYxbh5lNx5wYZE; wire [14:0] sIVqloL9MjkDXMyZqNgFi; wire [28:0] R5FT4wZn7DjE5FtgHFUm3E; wire [27:0] on0J0v1C0T4Vx5BAyNciCG; reg [31:0] zjMYjjAxK45sdDEQ0XFXOG; wire [27:0] xbDZHFjT9czSWoXqDrDalH; wire rIIATJviRgNIQoJq8fW3iH; wire [13:0] fWYsiC8varEjDaABQEOnHD; reg [13:0] jWzhv1CNrrkZ90yAhAoazF; wire [27:0] m6rhgeyCXShlzRN5AMh18G; wire [27:0] GJygrD3xsfw2DPQ22BhMnF; reg [27:0] rqeR6AxGoUnIpcf8RFZE0C; wire [29:0] uxJF4VESfR9zjMeGYtrIS; wire [15:0] a9YNARWK4HMkgu5zeMeFqB; wire [30:0] OJCxI8u48szx5fkdxbfWjF; wire [29:0] Nqy6crAgfKalgWwdaoPgWF; reg [31:0] UVyVvhhWLxLhiHSNKkfKfE; wire [29:0] VPMmTC28HmTVgoT6ZLk0CD; wire T4LoOhTfaEIFoiHehRN8gB; wire [14:0] z7KS1tRTiUNV07mMLJEuKG; reg [14:0] TKE1ENeioNod9UMhIzVfSH; wire [29:0] nkdnEk7YtJ3W7AmLNPDo; wire [29:0] y5KCvh2zjCyG1LFiVsUMYcD; reg [29:0] cZ0D6qUE7QWbwvVcyFlvNC; wire [31:0] zD10HQPaWNtGjDTMJz3GSH; wire [16:0] d9bLW3agjcpEpWrolrVdsmC; wire [32:0] QJOFvqfWKUFnEFOqoOrxWG; wire [31:0] z1qYldk164H9FNaPWpn6hF; reg [31:0] m47DvfSzOdN9OKy9YulLguB; wire cpmy5PzhVLGXdDoyCkUWiD; wire [15:0] LPQDAvbrOjkrOtmk9vzPJB; reg [15:0] agalUIcyHoMvnBXt7uR1FE; reg [15:0] VDuk3ojf4kqPZHi2nVzzSD [0:1]; wire [15:0] xzmEHvAakc16M7C3TuYQlF [0:1]; wire [15:0] n6vRpiFqkFIHzpDYbJGYiD; wire [15:0] q3w3Ce5AlDM2h7wxTsVajWB; wire XWhO1jBhWS8epPquTZyFzG; assign d2oEus6jJ0McV6ih95Y1AG = h4h0SDZC9CQgXKPbimISL3; assign Y8nU1xjYWVI5dgYrgIlsCE = d2oEus6jJ0McV6ih95Y1AG[31:30]; assign igWwj37zoLbvMLlrefWxbF = 2'b01 <= Y8nU1xjYWVI5dgYrgIlsCE; assign PtqvgNqZpdLWxF206ad9XC = (igWwj37zoLbvMLlrefWxbF == 1'b0 ? 1'b0 : 1'b1); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : c5cs351kKqE0paJffH20ksB if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin Td50TMNbpGWZYlXbqSVvTG <= 1'b0; end else begin Td50TMNbpGWZYlXbqSVvTG <= PtqvgNqZpdLWxF206ad9XC; end end assign f57E5i0241V1QEgB58U5YC = (igWwj37zoLbvMLlrefWxbF == 1'b0 ? 2'b00 : 2'b01); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : HfJzyVbuSarQZwy9cyUpkF if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin htY8XTFJI2P1kmv6r9UdwG <= 2'b00; end else begin htY8XTFJI2P1kmv6r9UdwG <= f57E5i0241V1QEgB58U5YC; end end assign mAB2T9yHc4paNxEah9oqhC = {htY8XTFJI2P1kmv6r9UdwG, 2'b01}; assign KhlHtRMHix8XvnicPL5XdC = {Td50TMNbpGWZYlXbqSVvTG, 2'b00}; assign lFIFc1FMCEhdqlYwYW5oSD = ({1'b0, mAB2T9yHc4paNxEah9oqhC}) + ({2'b0, KhlHtRMHix8XvnicPL5XdC}); assign OP66o1rkZm1IVPqs42DN1C = (lFIFc1FMCEhdqlYwYW5oSD[4] != 1'b0 ? 4'b1111 : lFIFc1FMCEhdqlYwYW5oSD[3:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : g2Pn1ppBtUFLbR5PDvbUBWE if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin p9JdL74lJmHuomPqcevLHkB <= 32'b00000000000000000000000000000000; end else begin p9JdL74lJmHuomPqcevLHkB <= d2oEus6jJ0McV6ih95Y1AG; end end assign RraIPFfLtZsHXCwvliBhwH = p9JdL74lJmHuomPqcevLHkB[31:28]; assign X1dRLKXI3e3fN1rBDqxex = OP66o1rkZm1IVPqs42DN1C <= RraIPFfLtZsHXCwvliBhwH; assign WN8EiF2jALV8OH7W7KXXaG = {Td50TMNbpGWZYlXbqSVvTG, X1dRLKXI3e3fN1rBDqxex}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : x0pPRCM2OL5qJQN0lZwEoL if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin OAnPRhXN1f3PXR2YrHATCE <= 2'b00; end else begin OAnPRhXN1f3PXR2YrHATCE <= WN8EiF2jALV8OH7W7KXXaG; end end assign bj4j66oAvfSpNoFLxGto1G = {htY8XTFJI2P1kmv6r9UdwG, 2'b00}; assign jZJyU4ZP4ChZ5K7R8RriDE = (X1dRLKXI3e3fN1rBDqxex == 1'b0 ? bj4j66oAvfSpNoFLxGto1G : OP66o1rkZm1IVPqs42DN1C); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : WwUtsWIaw94Jy54QEMHzF if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin aIuu8srO6WIrizhN08OyGG <= 4'b0000; end else begin aIuu8srO6WIrizhN08OyGG <= jZJyU4ZP4ChZ5K7R8RriDE; end end assign la6NpbM3xhaAGZJpg3nLdG = {aIuu8srO6WIrizhN08OyGG, 2'b01}; assign UAlS8hgEMaTiqrIEBR7P8D = {OAnPRhXN1f3PXR2YrHATCE, 2'b00}; assign DB14wLF62mIfBaTI6vec6B = ({1'b0, la6NpbM3xhaAGZJpg3nLdG}) + ({3'b0, UAlS8hgEMaTiqrIEBR7P8D}); assign Uf33riUqPe3QbDaMY9cxIE = (DB14wLF62mIfBaTI6vec6B[6] != 1'b0 ? 6'b111111 : DB14wLF62mIfBaTI6vec6B[5:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : YSqZgetA5RNmyz8MPSmuEG if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin EVGDcYjDYMyphmfUWLd40D <= 32'b00000000000000000000000000000000; end else begin EVGDcYjDYMyphmfUWLd40D <= p9JdL74lJmHuomPqcevLHkB; end end assign Ir5J1cq3X4AtmuV2rRCWJE = EVGDcYjDYMyphmfUWLd40D[31:26]; assign IfNgpXh3L8PgtuQ9riD96F = Uf33riUqPe3QbDaMY9cxIE <= Ir5J1cq3X4AtmuV2rRCWJE; assign rjTlAhUbkx4xhnY4CEQzSE = {OAnPRhXN1f3PXR2YrHATCE, IfNgpXh3L8PgtuQ9riD96F}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : DgFbJwbmEnKI37yyqDcNIG if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin Bb4Fv4CfcqYV9v1KrOFClE <= 3'b000; end else begin Bb4Fv4CfcqYV9v1KrOFClE <= rjTlAhUbkx4xhnY4CEQzSE; end end assign QBdSjsMcWKRY5gwAzbQLsH = {aIuu8srO6WIrizhN08OyGG, 2'b00}; assign SxeI6Ebz4W3cAlBHX6N7HE = (IfNgpXh3L8PgtuQ9riD96F == 1'b0 ? QBdSjsMcWKRY5gwAzbQLsH : Uf33riUqPe3QbDaMY9cxIE); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : aNYj5lvbs8Fnxy53OXvirH if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin a8prI6r0sJOb3uF5oZRDzvE <= 6'b000000; end else begin a8prI6r0sJOb3uF5oZRDzvE <= SxeI6Ebz4W3cAlBHX6N7HE; end end assign f4gekvhdG5D2vtDRQuIsRWD = {a8prI6r0sJOb3uF5oZRDzvE, 2'b01}; assign HlCg528B0DhdId48qwIzID = {Bb4Fv4CfcqYV9v1KrOFClE, 2'b00}; assign DdWFbmNZw3i61r2Flc3lJG = ({1'b0, f4gekvhdG5D2vtDRQuIsRWD}) + ({4'b0, HlCg528B0DhdId48qwIzID}); assign C1ig1Tdqfa5ultBNsDcUCH = (DdWFbmNZw3i61r2Flc3lJG[8] != 1'b0 ? 8'b11111111 : DdWFbmNZw3i61r2Flc3lJG[7:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : o0HUgiqSTXgxerKYJHQpdoH if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin RRY6uI32JPF7cgRt2ALKpD <= 32'b00000000000000000000000000000000; end else begin RRY6uI32JPF7cgRt2ALKpD <= EVGDcYjDYMyphmfUWLd40D; end end assign gMvZmbcqZ0DqgJ5sO7TczG = RRY6uI32JPF7cgRt2ALKpD[31:24]; assign WPfmCIzxCRH3PoV577VFZ = C1ig1Tdqfa5ultBNsDcUCH <= gMvZmbcqZ0DqgJ5sO7TczG; assign mIsPzyrzh6zMIEjXAztfSH = {Bb4Fv4CfcqYV9v1KrOFClE, WPfmCIzxCRH3PoV577VFZ}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : r8CDQXfJLKAhqXMOxSnRJE if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin W6W5MbHcLxMQiocqir3EcD <= 4'b0000; end else begin W6W5MbHcLxMQiocqir3EcD <= mIsPzyrzh6zMIEjXAztfSH; end end assign b6B3OCDRqPO9Qa8fvVfkrL = {a8prI6r0sJOb3uF5oZRDzvE, 2'b00}; assign c0V0PWcNTcAtWfHHZo9oCB = (WPfmCIzxCRH3PoV577VFZ == 1'b0 ? b6B3OCDRqPO9Qa8fvVfkrL : C1ig1Tdqfa5ultBNsDcUCH); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : TK10f4FbeDHxD5MzedXqjE if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin fCoWIZZx9VblaWmYgt13x <= 8'b00000000; end else begin fCoWIZZx9VblaWmYgt13x <= c0V0PWcNTcAtWfHHZo9oCB; end end assign btCYaoeB2JmWOR056EcY2C = {fCoWIZZx9VblaWmYgt13x, 2'b01}; assign IgY2MGVmpmzbfdJvodzhYH = {W6W5MbHcLxMQiocqir3EcD, 2'b00}; assign x2qOSwxaMdgo7eci0FxvvcF = ({1'b0, btCYaoeB2JmWOR056EcY2C}) + ({5'b0, IgY2MGVmpmzbfdJvodzhYH}); assign baKrdskhfkPzPlkAHW54rF = (x2qOSwxaMdgo7eci0FxvvcF[10] != 1'b0 ? 10'b1111111111 : x2qOSwxaMdgo7eci0FxvvcF[9:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : T84SIUDYmHxjd2ywg6pY9 if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin JnW70VzeuX4yEHMB8XIxSE <= 32'b00000000000000000000000000000000; end else begin JnW70VzeuX4yEHMB8XIxSE <= RRY6uI32JPF7cgRt2ALKpD; end end assign p3SL7wYX8SBQnC0oYVuIuHF = JnW70VzeuX4yEHMB8XIxSE[31:22]; assign q48UwMWOiN7vMKVlbAH62tG = baKrdskhfkPzPlkAHW54rF <= p3SL7wYX8SBQnC0oYVuIuHF; assign xTGR6ce6S4BzV4dkYyod4F = {W6W5MbHcLxMQiocqir3EcD, q48UwMWOiN7vMKVlbAH62tG}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : eqqkIKQHHL0nSk056vyEfF if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin jXOqwspdsCISwsGhcWqtUE <= 5'b00000; end else begin jXOqwspdsCISwsGhcWqtUE <= xTGR6ce6S4BzV4dkYyod4F; end end assign fkhBlawaiECm3AKyJOvEc = {fCoWIZZx9VblaWmYgt13x, 2'b00}; assign QDLMg0wJNF3uVvsVP11Se = (q48UwMWOiN7vMKVlbAH62tG == 1'b0 ? fkhBlawaiECm3AKyJOvEc : baKrdskhfkPzPlkAHW54rF); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : ta6nlbGoEbbBQly2tMoP5C if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin kfyELMjsnnzaUx6iYLK1a <= 10'b0000000000; end else begin kfyELMjsnnzaUx6iYLK1a <= QDLMg0wJNF3uVvsVP11Se; end end assign j3mLQ1yo2zmp8dnGzKOW5qB = {kfyELMjsnnzaUx6iYLK1a, 2'b01}; assign H5Q1sQZfYTS1fDeRqymzvG = {jXOqwspdsCISwsGhcWqtUE, 2'b00}; assign i7x1l0whvlbCztZ8yv9iwE = ({1'b0, j3mLQ1yo2zmp8dnGzKOW5qB}) + ({6'b0, H5Q1sQZfYTS1fDeRqymzvG}); assign ztLkXaVGX3w4pEn1xeRqMC = (i7x1l0whvlbCztZ8yv9iwE[12] != 1'b0 ? 12'b111111111111 : i7x1l0whvlbCztZ8yv9iwE[11:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : r6S7UYwuR8Ixw8Lmwe9W8KE if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin rMhu2oApltCVSYS5itmY0C <= 32'b00000000000000000000000000000000; end else begin rMhu2oApltCVSYS5itmY0C <= JnW70VzeuX4yEHMB8XIxSE; end end assign r46CEAiCE4Ch2WNWkeHtNeF = rMhu2oApltCVSYS5itmY0C[31:20]; assign PloSd07HvtUIeQYlow2DsD = ztLkXaVGX3w4pEn1xeRqMC <= r46CEAiCE4Ch2WNWkeHtNeF; assign wm9pXs3ggIACgFF4VQ65zG = {jXOqwspdsCISwsGhcWqtUE, PloSd07HvtUIeQYlow2DsD}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : x28YJ6sLjBQMYm398bLX0OC if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin YfPairRXLNNVGttdcC4jHC <= 6'b000000; end else begin YfPairRXLNNVGttdcC4jHC <= wm9pXs3ggIACgFF4VQ65zG; end end assign actzjOg0aKNbyOOWNABa6F = {kfyELMjsnnzaUx6iYLK1a, 2'b00}; assign l0kGuUM557NseEtaykZ1TID = (PloSd07HvtUIeQYlow2DsD == 1'b0 ? actzjOg0aKNbyOOWNABa6F : ztLkXaVGX3w4pEn1xeRqMC); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : Abpc1Ylh34fRxdRvHjZv7 if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin wBLoEXjrUx0g620zErfyIH <= 12'b000000000000; end else begin wBLoEXjrUx0g620zErfyIH <= l0kGuUM557NseEtaykZ1TID; end end assign jARRiz24LDX5CAkjjvpbMC = {wBLoEXjrUx0g620zErfyIH, 2'b01}; assign cOqqXZggK8lV63HuJIDU6C = {YfPairRXLNNVGttdcC4jHC, 2'b00}; assign g03PW5Zn8wGm996TsM3OlSG = ({1'b0, jARRiz24LDX5CAkjjvpbMC}) + ({7'b0, cOqqXZggK8lV63HuJIDU6C}); assign seXC0DlX19Qu2W9b6laBkF = (g03PW5Zn8wGm996TsM3OlSG[14] != 1'b0 ? 14'b11111111111111 : g03PW5Zn8wGm996TsM3OlSG[13:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : lvsMaaP5bWohwV7eCS6Ih if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin YuoRtO5uahqj9k1hlroeUD <= 32'b00000000000000000000000000000000; end else begin YuoRtO5uahqj9k1hlroeUD <= rMhu2oApltCVSYS5itmY0C; end end assign VJtd7Fl5sWCBbwZ7zVkiAH = YuoRtO5uahqj9k1hlroeUD[31:18]; assign DFiuspHBeirfq1ZvvofTRC = seXC0DlX19Qu2W9b6laBkF <= VJtd7Fl5sWCBbwZ7zVkiAH; assign ym9Sp6nhcDPOiwj0UyGXsC = {YfPairRXLNNVGttdcC4jHC, DFiuspHBeirfq1ZvvofTRC}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : A52ertO1i9dzNTTRoQFYZ if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin zQQJr5Rr8Ek603tPKykxHC <= 7'b0000000; end else begin zQQJr5Rr8Ek603tPKykxHC <= ym9Sp6nhcDPOiwj0UyGXsC; end end assign P1SxQfGkK55cR5k1YisfzE = {wBLoEXjrUx0g620zErfyIH, 2'b00}; assign tp0Xxl65VoHaM4O6FDb2N = (DFiuspHBeirfq1ZvvofTRC == 1'b0 ? P1SxQfGkK55cR5k1YisfzE : seXC0DlX19Qu2W9b6laBkF); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : r9aaNhIpaPxlclpq2W48eD if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin toUJwGxo7JfW2EzqeaegqD <= 14'b00000000000000; end else begin toUJwGxo7JfW2EzqeaegqD <= tp0Xxl65VoHaM4O6FDb2N; end end assign hqJrTgFxozMyPx7LnmLBzE = {toUJwGxo7JfW2EzqeaegqD, 2'b01}; assign i3H4mRdiwOgMnPaGpxPykE = {zQQJr5Rr8Ek603tPKykxHC, 2'b00}; assign IbH5QT2AXNs8KsoyD12ZfE = ({1'b0, hqJrTgFxozMyPx7LnmLBzE}) + ({8'b0, i3H4mRdiwOgMnPaGpxPykE}); assign V1kZ7bFxQFV1KrNlMFxWYG = (IbH5QT2AXNs8KsoyD12ZfE[16] != 1'b0 ? 16'b1111111111111111 : IbH5QT2AXNs8KsoyD12ZfE[15:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : UB4F966VLLxkmGZ0IGY51G if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin vAj4ixajCquQJTqGQyxOnB <= 32'b00000000000000000000000000000000; end else begin vAj4ixajCquQJTqGQyxOnB <= YuoRtO5uahqj9k1hlroeUD; end end assign O219BqtpHO98GKSgKS8BpE = vAj4ixajCquQJTqGQyxOnB[31:16]; assign FTmP9v6IJWTPVZpRmGRtIF = V1kZ7bFxQFV1KrNlMFxWYG <= O219BqtpHO98GKSgKS8BpE; assign pv1WByjbGdV1OSiqH0ksnC = {zQQJr5Rr8Ek603tPKykxHC, FTmP9v6IJWTPVZpRmGRtIF}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : c7pLAVb4q0zp9SmImNpMy5F if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin DfmgsE3iMkzCsirhmlRDSH <= 8'b00000000; end else begin DfmgsE3iMkzCsirhmlRDSH <= pv1WByjbGdV1OSiqH0ksnC; end end assign x40VeLX7J3a3tphEEkOgR2D = {toUJwGxo7JfW2EzqeaegqD, 2'b00}; assign n6crFALdZyJcOXZ3tAFGjWE = (FTmP9v6IJWTPVZpRmGRtIF == 1'b0 ? x40VeLX7J3a3tphEEkOgR2D : V1kZ7bFxQFV1KrNlMFxWYG); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : TmD5lx10ao7OSow20n40KH if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin q72w2glJ0iF1fL3kkboMy5C <= 16'b0000000000000000; end else begin q72w2glJ0iF1fL3kkboMy5C <= n6crFALdZyJcOXZ3tAFGjWE; end end assign eUkkETd043d2fZQk8jDNbG = {q72w2glJ0iF1fL3kkboMy5C, 2'b01}; assign ctWCGk8tDhNhqjRiNbiT8G = {DfmgsE3iMkzCsirhmlRDSH, 2'b00}; assign jtIl02WJwApYjH6zHw0ps = ({1'b0, eUkkETd043d2fZQk8jDNbG}) + ({9'b0, ctWCGk8tDhNhqjRiNbiT8G}); assign aEmD7oGZhl9CNV3Ln3b9jD = (jtIl02WJwApYjH6zHw0ps[18] != 1'b0 ? 18'b111111111111111111 : jtIl02WJwApYjH6zHw0ps[17:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : l3fzdqpAByu1sqIOkQhtH3F if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin u2ZdQtNDigVBNNBtq7C1PFC <= 32'b00000000000000000000000000000000; end else begin u2ZdQtNDigVBNNBtq7C1PFC <= vAj4ixajCquQJTqGQyxOnB; end end assign xUhkT9IaYCKujHljsYB4WB = u2ZdQtNDigVBNNBtq7C1PFC[31:14]; assign aEXdj8byA7uSgyb9LhSHuH = aEmD7oGZhl9CNV3Ln3b9jD <= xUhkT9IaYCKujHljsYB4WB; assign Yw6DjbSH20VSb4AH6J2ZW = {DfmgsE3iMkzCsirhmlRDSH, aEXdj8byA7uSgyb9LhSHuH}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : NLDk95Gtp0Xpqh8HvNrDKC if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin VlHUymZGBDkWniRKHnXeoE <= 9'b000000000; end else begin VlHUymZGBDkWniRKHnXeoE <= Yw6DjbSH20VSb4AH6J2ZW; end end assign BmC7Waj3h156ApBRR8vBkB = {q72w2glJ0iF1fL3kkboMy5C, 2'b00}; assign e6y0zTjYMJQBzfcOI5kwLeC = (aEXdj8byA7uSgyb9LhSHuH == 1'b0 ? BmC7Waj3h156ApBRR8vBkB : aEmD7oGZhl9CNV3Ln3b9jD); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : THTy90hfyvYqXVkE8CcRgG if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin goHRzycDTV9MFT2FCIUeIF <= 18'b000000000000000000; end else begin goHRzycDTV9MFT2FCIUeIF <= e6y0zTjYMJQBzfcOI5kwLeC; end end assign QLgRzXPFcx5iBqm0rMhzn = {goHRzycDTV9MFT2FCIUeIF, 2'b01}; assign xbtGwTj2py2rKQx3DwaqsH = {VlHUymZGBDkWniRKHnXeoE, 2'b00}; assign l5Svt4GkcCOLXXQwBiRIcD = ({1'b0, QLgRzXPFcx5iBqm0rMhzn}) + ({10'b0, xbtGwTj2py2rKQx3DwaqsH}); assign wCUr9vYed0L827ZSFIusEB = (l5Svt4GkcCOLXXQwBiRIcD[20] != 1'b0 ? 20'b11111111111111111111 : l5Svt4GkcCOLXXQwBiRIcD[19:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : Wi3GKYc8qmHzWSUSCWfLqC if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin yI0NKYDzTZw44KqJ9a3zC <= 32'b00000000000000000000000000000000; end else begin yI0NKYDzTZw44KqJ9a3zC <= u2ZdQtNDigVBNNBtq7C1PFC; end end assign bkWNTMVtSZYFA4nZXmoiEG = yI0NKYDzTZw44KqJ9a3zC[31:12]; assign vlYCGljOoPPGkfFDbGHWcC = wCUr9vYed0L827ZSFIusEB <= bkWNTMVtSZYFA4nZXmoiEG; assign SZm8Zt2WiFh8VGkrN5GsuC = {VlHUymZGBDkWniRKHnXeoE, vlYCGljOoPPGkfFDbGHWcC}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : lHhT3gqQkx9RTwHwtL7LeC if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin e56HDsGesAEqHwWeqzouMF <= 10'b0000000000; end else begin e56HDsGesAEqHwWeqzouMF <= SZm8Zt2WiFh8VGkrN5GsuC; end end assign zLl2QCAAjWMixlTOkaGHiE = {goHRzycDTV9MFT2FCIUeIF, 2'b00}; assign PcExrzPwT7phvvgF45pQHH = (vlYCGljOoPPGkfFDbGHWcC == 1'b0 ? zLl2QCAAjWMixlTOkaGHiE : wCUr9vYed0L827ZSFIusEB); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : i9eBCUMqIE3L7n0V9baxa2F if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin Wz90RhDyGBtEdtGrJ0VTZF <= 20'b00000000000000000000; end else begin Wz90RhDyGBtEdtGrJ0VTZF <= PcExrzPwT7phvvgF45pQHH; end end assign s2ByO9sLopwaaKB3OlviZB = {Wz90RhDyGBtEdtGrJ0VTZF, 2'b01}; assign SRZlivglW4iODt3ZWa6YAB = {e56HDsGesAEqHwWeqzouMF, 2'b00}; assign mTVvj9euDcz3QKkAdcmZOD = ({1'b0, s2ByO9sLopwaaKB3OlviZB}) + ({11'b0, SRZlivglW4iODt3ZWa6YAB}); assign ay59snlUFLNfqFr9K8OyMB = (mTVvj9euDcz3QKkAdcmZOD[22] != 1'b0 ? 22'b1111111111111111111111 : mTVvj9euDcz3QKkAdcmZOD[21:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : JxAPLal5Cdfhkgjtyzw9d if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin VrDvujAzBpk1JUnt3i3jrD <= 32'b00000000000000000000000000000000; end else begin VrDvujAzBpk1JUnt3i3jrD <= yI0NKYDzTZw44KqJ9a3zC; end end assign nXG6pKWoysTLlamoZb1kUC = VrDvujAzBpk1JUnt3i3jrD[31:10]; assign FVZq6SQWJqDew38uj3ZwuF = ay59snlUFLNfqFr9K8OyMB <= nXG6pKWoysTLlamoZb1kUC; assign UJGgN0K4zoVMt8OzpDRhbB = {e56HDsGesAEqHwWeqzouMF, FVZq6SQWJqDew38uj3ZwuF}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : GxjkjjAOj44SCVWlUX1tY if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin ElZOyt1VjSkVNH6qpuxaXG <= 11'b00000000000; end else begin ElZOyt1VjSkVNH6qpuxaXG <= UJGgN0K4zoVMt8OzpDRhbB; end end assign w0u8eyeEsFecynkh04cF1lC = {Wz90RhDyGBtEdtGrJ0VTZF, 2'b00}; assign WXHkYoAaBaLUFbVOCc8VxD = (FVZq6SQWJqDew38uj3ZwuF == 1'b0 ? w0u8eyeEsFecynkh04cF1lC : ay59snlUFLNfqFr9K8OyMB); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : d6h65HOwLiX9kWQsaGF4qnC if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin pNjnAf3CRLybq0T318tpZB <= 22'b0000000000000000000000; end else begin pNjnAf3CRLybq0T318tpZB <= WXHkYoAaBaLUFbVOCc8VxD; end end assign pUZF40VeZ6xEJvpR7Es8FG = {pNjnAf3CRLybq0T318tpZB, 2'b01}; assign CZy9D9fjHBHcfkgtp0KTFH = {ElZOyt1VjSkVNH6qpuxaXG, 2'b00}; assign kLW7ETLJg3f0fhJvPfzamC = ({1'b0, pUZF40VeZ6xEJvpR7Es8FG}) + ({12'b0, CZy9D9fjHBHcfkgtp0KTFH}); assign jV8kLyXAcS3FCyqURyzmO = (kLW7ETLJg3f0fhJvPfzamC[24] != 1'b0 ? 24'b111111111111111111111111 : kLW7ETLJg3f0fhJvPfzamC[23:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : KFx91owMzgsCl6NpENL6wF if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin iLdfuowoyk1MtRrU15MG4C <= 32'b00000000000000000000000000000000; end else begin iLdfuowoyk1MtRrU15MG4C <= VrDvujAzBpk1JUnt3i3jrD; end end assign q9f5spD683cNlZnQf56m4ZE = iLdfuowoyk1MtRrU15MG4C[31:8]; assign qE7EncjwDfib2QclnYwSgG = jV8kLyXAcS3FCyqURyzmO <= q9f5spD683cNlZnQf56m4ZE; assign PPmIvwimSHZwNXz56Jo5FF = {ElZOyt1VjSkVNH6qpuxaXG, qE7EncjwDfib2QclnYwSgG}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : mlbpF5PDgS6CPvuh9fETwH if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin s7H3AIDyv88anihczWgA1F <= 12'b000000000000; end else begin s7H3AIDyv88anihczWgA1F <= PPmIvwimSHZwNXz56Jo5FF; end end assign fjwwR4v4yEuDBPgyT1rTBE = {pNjnAf3CRLybq0T318tpZB, 2'b00}; assign JRbiQknn0l3SAzJguSaDIE = (qE7EncjwDfib2QclnYwSgG == 1'b0 ? fjwwR4v4yEuDBPgyT1rTBE : jV8kLyXAcS3FCyqURyzmO); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : wCPDI5egX7bGmr1qgDF9WE if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin ebaB1Kw2OvZfbCMRd7RH4G <= 24'b000000000000000000000000; end else begin ebaB1Kw2OvZfbCMRd7RH4G <= JRbiQknn0l3SAzJguSaDIE; end end assign WOq3F3uShD744l8tfCN3PC = {ebaB1Kw2OvZfbCMRd7RH4G, 2'b01}; assign te9YCAmyrsrdkIOdNQ10YB = {s7H3AIDyv88anihczWgA1F, 2'b00}; assign r0mlnEduB1ta4alefYkcSzF = ({1'b0, WOq3F3uShD744l8tfCN3PC}) + ({13'b0, te9YCAmyrsrdkIOdNQ10YB}); assign chc7OKgA3bugXJCo3yas7F = (r0mlnEduB1ta4alefYkcSzF[26] != 1'b0 ? 26'b11111111111111111111111111 : r0mlnEduB1ta4alefYkcSzF[25:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : lAj0wFX3ymFHEKGROpovNF if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin lEZvI5hvOIId49rKN6EG9B <= 32'b00000000000000000000000000000000; end else begin lEZvI5hvOIId49rKN6EG9B <= iLdfuowoyk1MtRrU15MG4C; end end assign d4IpN7AeFzlW8PIZDtHBNhH = lEZvI5hvOIId49rKN6EG9B[31:6]; assign kdK0vZeghYKX1pPI7TOLUG = chc7OKgA3bugXJCo3yas7F <= d4IpN7AeFzlW8PIZDtHBNhH; assign vIkIEBTGTAhgY525Xqzf1E = {s7H3AIDyv88anihczWgA1F, kdK0vZeghYKX1pPI7TOLUG}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : RTZmiZqqJJb7QmO7j7Q28E if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin Igu3qoayK7OqaCOGUvR5mH <= 13'b0000000000000; end else begin Igu3qoayK7OqaCOGUvR5mH <= vIkIEBTGTAhgY525Xqzf1E; end end assign uR89cXy8xlRQIE7YbWSVVF = {ebaB1Kw2OvZfbCMRd7RH4G, 2'b00}; assign jWK6QZgHeyt3ftPSKbIyaD = (kdK0vZeghYKX1pPI7TOLUG == 1'b0 ? uR89cXy8xlRQIE7YbWSVVF : chc7OKgA3bugXJCo3yas7F); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : b65fXEthqOsaOZSgRWDuCE if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin I9gVg5rOTUbEKRzS4CERmD <= 26'b00000000000000000000000000; end else begin I9gVg5rOTUbEKRzS4CERmD <= jWK6QZgHeyt3ftPSKbIyaD; end end assign UTCgRY29pVn3brpE5SMH2C = {I9gVg5rOTUbEKRzS4CERmD, 2'b01}; assign v43le787IqXWHekLEH8sc1F = {Igu3qoayK7OqaCOGUvR5mH, 2'b00}; assign ERrwsqMxpQKfcAVllHsC = ({1'b0, UTCgRY29pVn3brpE5SMH2C}) + ({14'b0, v43le787IqXWHekLEH8sc1F}); assign NztI2AQnSAdBX3RAcWFzi = (ERrwsqMxpQKfcAVllHsC[28] != 1'b0 ? 28'b1111111111111111111111111111 : ERrwsqMxpQKfcAVllHsC[27:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : zZfAZ5rDiGQaCF1bs2ULU if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin nY5HJQdvwbdw1Z09MGQJdD <= 32'b00000000000000000000000000000000; end else begin nY5HJQdvwbdw1Z09MGQJdD <= lEZvI5hvOIId49rKN6EG9B; end end assign ZH59np0e4GT0PI42ZDK96D = nY5HJQdvwbdw1Z09MGQJdD[31:4]; assign qvx4HYpxmuqVBKosKL9nDF = NztI2AQnSAdBX3RAcWFzi <= ZH59np0e4GT0PI42ZDK96D; assign vXQqwFz0Mq5pyOl5hUGpTE = {Igu3qoayK7OqaCOGUvR5mH, qvx4HYpxmuqVBKosKL9nDF}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : Ns4fsEtlsMtY3wmIYgUi9D if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin XSv77atgil9CALLij3LDU <= 14'b00000000000000; end else begin XSv77atgil9CALLij3LDU <= vXQqwFz0Mq5pyOl5hUGpTE; end end assign fqeYT46R9tLTDvWKi4sZDC = {I9gVg5rOTUbEKRzS4CERmD, 2'b00}; assign FQVTrSjADBrb3DyvHSAwpC = (qvx4HYpxmuqVBKosKL9nDF == 1'b0 ? fqeYT46R9tLTDvWKi4sZDC : NztI2AQnSAdBX3RAcWFzi); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : m22lc0RW2bbIMYyadLgFhD if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin k2Wyo4gBkJTLcHbPeag55GC <= 28'b0000000000000000000000000000; end else begin k2Wyo4gBkJTLcHbPeag55GC <= FQVTrSjADBrb3DyvHSAwpC; end end assign bb45jO7OrRC3XbD8zJ6puE = {k2Wyo4gBkJTLcHbPeag55GC, 2'b01}; assign XXiXbfRxJuy8atUhokFqtC = {XSv77atgil9CALLij3LDU, 2'b00}; assign UW4b3bm76Bs6tI3IYkPZIE = ({1'b0, bb45jO7OrRC3XbD8zJ6puE}) + ({15'b0, XXiXbfRxJuy8atUhokFqtC}); assign q55ENw2wkQaVRklvIu1LrF = (UW4b3bm76Bs6tI3IYkPZIE[30] != 1'b0 ? 30'b111111111111111111111111111111 : UW4b3bm76Bs6tI3IYkPZIE[29:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : s9xKMW8bbefctNY9iigvNBC if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin aJrV9N3G9wp8U0g9mfcyX <= 32'b00000000000000000000000000000000; end else begin aJrV9N3G9wp8U0g9mfcyX <= nY5HJQdvwbdw1Z09MGQJdD; end end assign ZYrtxtrqxr2hmg5PKUYcOG = aJrV9N3G9wp8U0g9mfcyX[31:2]; assign X1QJVAhYCy1C1RlcRQ7ehC = q55ENw2wkQaVRklvIu1LrF <= ZYrtxtrqxr2hmg5PKUYcOG; assign cLzalZ4N3AQH17rH3HxvHG = {XSv77atgil9CALLij3LDU, X1QJVAhYCy1C1RlcRQ7ehC}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : oDLsLJn2kyFBG6g0aa6kxD if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin FoKnmJHxBvoWITgnEM5uGB <= 15'b000000000000000; end else begin FoKnmJHxBvoWITgnEM5uGB <= cLzalZ4N3AQH17rH3HxvHG; end end assign u4MPAwPCLIAgQPn96oG4E2C = {k2Wyo4gBkJTLcHbPeag55GC, 2'b00}; assign muL6drwYusIoOSLLD6cQME = (X1QJVAhYCy1C1RlcRQ7ehC == 1'b0 ? u4MPAwPCLIAgQPn96oG4E2C : q55ENw2wkQaVRklvIu1LrF); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : r4wvZUUnsyepUkKB0zo9yF if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin ECSbb2HpHz8MkgOToIfkRB <= 30'b000000000000000000000000000000; end else begin ECSbb2HpHz8MkgOToIfkRB <= muL6drwYusIoOSLLD6cQME; end end assign pUbtxeEGlqbH77tEidOseF = {ECSbb2HpHz8MkgOToIfkRB, 2'b01}; assign OBIn9RfqwS76ifr6ctbJcC = {FoKnmJHxBvoWITgnEM5uGB, 2'b00}; assign Vd09OCdvDhHzYbNi8eFYqD = ({1'b0, pUbtxeEGlqbH77tEidOseF}) + ({16'b0, OBIn9RfqwS76ifr6ctbJcC}); assign x9dWBNZVozdT9sZOUOShSwE = (Vd09OCdvDhHzYbNi8eFYqD[32] != 1'b0 ? 32'b11111111111111111111111111111111 : Vd09OCdvDhHzYbNi8eFYqD[31:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : b7HQI8ZyJUamitTLsYSRYD if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin c1Fi1DCmwETWogyXFP0luXH <= 32'b00000000000000000000000000000000; end else begin c1Fi1DCmwETWogyXFP0luXH <= aJrV9N3G9wp8U0g9mfcyX; end end assign BQlKwJMG1iIAM1sM8WOwZD = x9dWBNZVozdT9sZOUOShSwE <= c1Fi1DCmwETWogyXFP0luXH; assign U6NVSwrrDlIXWmZMGhGnGF = {FoKnmJHxBvoWITgnEM5uGB, BQlKwJMG1iIAM1sM8WOwZD}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : PQ6Dxe1LpWhxaMX4UzuP1C if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin CNCrh0XltTO38hUhsOK89E <= 16'b0000000000000000; end else begin CNCrh0XltTO38hUhsOK89E <= U6NVSwrrDlIXWmZMGhGnGF; end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : UwIvVC5FAB8rbKWhh44Rd if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin tuyMU89x2cRtnHZbS629ED[0] <= 16'b0000000000000000; tuyMU89x2cRtnHZbS629ED[1] <= 16'b0000000000000000; end else begin tuyMU89x2cRtnHZbS629ED[0] <= X4jT0JtvhLt1PtInljBofC[0]; tuyMU89x2cRtnHZbS629ED[1] <= X4jT0JtvhLt1PtInljBofC[1]; end end assign FTPlQQTDuHArhica0zG5YE = tuyMU89x2cRtnHZbS629ED[1]; assign X4jT0JtvhLt1PtInljBofC[0] = CNCrh0XltTO38hUhsOK89E; assign X4jT0JtvhLt1PtInljBofC[1] = tuyMU89x2cRtnHZbS629ED[0]; assign ztGXs97JmxTgacz6ch5gZB = FTPlQQTDuHArhica0zG5YE; assign j71O4t3Nm1w5MRqcbOUNtHF = ztGXs97JmxTgacz6ch5gZB; assign kilI6xSQxSJzoqPMjerk6G = b0pPxQrhAhYENzTiTGGny5G; assign FbKbMjw44CL9zGZx7WXzGF = kilI6xSQxSJzoqPMjerk6G[31:30]; assign fB6UnuVq9iLH8XGHOxxXZD = 2'b01 <= FbKbMjw44CL9zGZx7WXzGF; assign UPTJ0KHCAkQKe7namSEKjC = (fB6UnuVq9iLH8XGHOxxXZD == 1'b0 ? 1'b0 : 1'b1); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : q7kpFFSAp3c8yXq18kqRPlH if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin YWY1tbo2DIf9KVzn8BwzCG <= 1'b0; end else begin YWY1tbo2DIf9KVzn8BwzCG <= UPTJ0KHCAkQKe7namSEKjC; end end assign z1nwdQwUNbMUELLx9AUfwkH = (fB6UnuVq9iLH8XGHOxxXZD == 1'b0 ? 2'b00 : 2'b01); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : mGxjPCgfoJVG8VaVTi6nAD if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin MEBenkOBGLeR7FTQrrn3MD <= 2'b00; end else begin MEBenkOBGLeR7FTQrrn3MD <= z1nwdQwUNbMUELLx9AUfwkH; end end assign O6EltwTicLhBoBnh9C7QlF = {MEBenkOBGLeR7FTQrrn3MD, 2'b01}; assign WDqWbhmj05r4Wjj5vIY3CE = {YWY1tbo2DIf9KVzn8BwzCG, 2'b00}; assign cxg6xJXOtsYvHf3YKjaqmH = ({1'b0, O6EltwTicLhBoBnh9C7QlF}) + ({2'b0, WDqWbhmj05r4Wjj5vIY3CE}); assign vzZzLR6yNvm5R3q77DDCBG = (cxg6xJXOtsYvHf3YKjaqmH[4] != 1'b0 ? 4'b1111 : cxg6xJXOtsYvHf3YKjaqmH[3:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : AkZmervM1XCNmAMWEX2SNF if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin ecTpLKJNtox43CqRvB7TqH <= 32'b00000000000000000000000000000000; end else begin ecTpLKJNtox43CqRvB7TqH <= kilI6xSQxSJzoqPMjerk6G; end end assign YX0TWRD0dHUDqZu2WRc64C = ecTpLKJNtox43CqRvB7TqH[31:28]; assign FCe1MyFX72qFVD3Hy9hPUE = vzZzLR6yNvm5R3q77DDCBG <= YX0TWRD0dHUDqZu2WRc64C; assign j6CDlg9BLVqvfP3aItxlu6G = {YWY1tbo2DIf9KVzn8BwzCG, FCe1MyFX72qFVD3Hy9hPUE}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : o3RaoMv27VvD8Yv8OWRmMaC if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin wEKIGBrNcPO2iCCXrGUIu <= 2'b00; end else begin wEKIGBrNcPO2iCCXrGUIu <= j6CDlg9BLVqvfP3aItxlu6G; end end assign d3qzATGoyxtZcYJcgfDfbeH = {MEBenkOBGLeR7FTQrrn3MD, 2'b00}; assign nOloqK6lS4ZdzwyM1eUzUB = (FCe1MyFX72qFVD3Hy9hPUE == 1'b0 ? d3qzATGoyxtZcYJcgfDfbeH : vzZzLR6yNvm5R3q77DDCBG); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : rBKgJ3MbibC0sk8FQNg16C if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin wpq9P4PBi8CGLKpUN7fWZB <= 4'b0000; end else begin wpq9P4PBi8CGLKpUN7fWZB <= nOloqK6lS4ZdzwyM1eUzUB; end end assign o65FJTz0B7IXjYcgfpVqSZB = {wpq9P4PBi8CGLKpUN7fWZB, 2'b01}; assign C47tZ0C1xf5jlTyv6MLJdF = {wEKIGBrNcPO2iCCXrGUIu, 2'b00}; assign lzW16GgG5bSiyHby6MJi7F = ({1'b0, o65FJTz0B7IXjYcgfpVqSZB}) + ({3'b0, C47tZ0C1xf5jlTyv6MLJdF}); assign o8P0gThAuIs85SmAegMaBdC = (lzW16GgG5bSiyHby6MJi7F[6] != 1'b0 ? 6'b111111 : lzW16GgG5bSiyHby6MJi7F[5:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : mIh3pRwzFJZsKoQKGsZmjF if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin NKytYt7HRGpr10Je7y72bD <= 32'b00000000000000000000000000000000; end else begin NKytYt7HRGpr10Je7y72bD <= ecTpLKJNtox43CqRvB7TqH; end end assign r5YWTZbOV1ZMPt3R1VWQsEF = NKytYt7HRGpr10Je7y72bD[31:26]; assign claoCCs3pNDgkEZUVS4BEC = o8P0gThAuIs85SmAegMaBdC <= r5YWTZbOV1ZMPt3R1VWQsEF; assign QKjfaK9XJfQuzgSPqcdG = {wEKIGBrNcPO2iCCXrGUIu, claoCCs3pNDgkEZUVS4BEC}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : MgcwL6ZAx48Vsp1Fzaa7KB if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin PVfspm0nrz7RTrj71zZK2E <= 3'b000; end else begin PVfspm0nrz7RTrj71zZK2E <= QKjfaK9XJfQuzgSPqcdG; end end assign bcdChZWFB9riH389qHJhvE = {wpq9P4PBi8CGLKpUN7fWZB, 2'b00}; assign JT69Ak8v7evsLSjX2WQmM = (claoCCs3pNDgkEZUVS4BEC == 1'b0 ? bcdChZWFB9riH389qHJhvE : o8P0gThAuIs85SmAegMaBdC); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : TwbveR48UHNtsNtTRIcxoG if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin t9R7A1peR6CuzTzZAm3HwC <= 6'b000000; end else begin t9R7A1peR6CuzTzZAm3HwC <= JT69Ak8v7evsLSjX2WQmM; end end assign QOFovA9T9qIZcEqTAPhtOF = {t9R7A1peR6CuzTzZAm3HwC, 2'b01}; assign iar9KCTPqGuEmE9kiyh5vE = {PVfspm0nrz7RTrj71zZK2E, 2'b00}; assign gCZzU6M0PYvvj8GKTwHOiG = ({1'b0, QOFovA9T9qIZcEqTAPhtOF}) + ({4'b0, iar9KCTPqGuEmE9kiyh5vE}); assign f1zvQhGH1CAcbvWG7t74yHC = (gCZzU6M0PYvvj8GKTwHOiG[8] != 1'b0 ? 8'b11111111 : gCZzU6M0PYvvj8GKTwHOiG[7:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : l7lXbR7aM97AGYv5180gpKC if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin Z4I0KdM2JVi87xjTMS96pG <= 32'b00000000000000000000000000000000; end else begin Z4I0KdM2JVi87xjTMS96pG <= NKytYt7HRGpr10Je7y72bD; end end assign nvyG06fFyy1jvHC47zz9RB = Z4I0KdM2JVi87xjTMS96pG[31:24]; assign cHWq2LRdov1nvfvvjvk3TG = f1zvQhGH1CAcbvWG7t74yHC <= nvyG06fFyy1jvHC47zz9RB; assign l1XFmcvlNKvaQmQZV9JV9jF = {PVfspm0nrz7RTrj71zZK2E, cHWq2LRdov1nvfvvjvk3TG}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : h5C5bOrOVtB5lkifyAma8hG if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin EokQF3Q771FYsuXM046eTE <= 4'b0000; end else begin EokQF3Q771FYsuXM046eTE <= l1XFmcvlNKvaQmQZV9JV9jF; end end assign DFG5jHCJODhySug0Ml3hXC = {t9R7A1peR6CuzTzZAm3HwC, 2'b00}; assign nqmUVeMYCM820YVZt5ilzG = (cHWq2LRdov1nvfvvjvk3TG == 1'b0 ? DFG5jHCJODhySug0Ml3hXC : f1zvQhGH1CAcbvWG7t74yHC); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : wZt1rb1BWMOZfNVRu8MlsG if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin f0Pv94BMpwnCMzWcufXc6hF <= 8'b00000000; end else begin f0Pv94BMpwnCMzWcufXc6hF <= nqmUVeMYCM820YVZt5ilzG; end end assign KbzFknNUACxVWcnzlxJfPH = {f0Pv94BMpwnCMzWcufXc6hF, 2'b01}; assign vQdMrvqDo8qF2kLKQ7AeXC = {EokQF3Q771FYsuXM046eTE, 2'b00}; assign MmjkPa4HYQ1KxOVnGr5TS = ({1'b0, KbzFknNUACxVWcnzlxJfPH}) + ({5'b0, vQdMrvqDo8qF2kLKQ7AeXC}); assign KiJFVa7Kln3PVycUSEnQNG = (MmjkPa4HYQ1KxOVnGr5TS[10] != 1'b0 ? 10'b1111111111 : MmjkPa4HYQ1KxOVnGr5TS[9:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : I33DRI27ZVR2M7fm8YlLxG if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin npDxBmN6dOapdh7YCQNR6E <= 32'b00000000000000000000000000000000; end else begin npDxBmN6dOapdh7YCQNR6E <= Z4I0KdM2JVi87xjTMS96pG; end end assign l9uTQkxnOKF0VsYALlWDi = npDxBmN6dOapdh7YCQNR6E[31:22]; assign df9yw7V8ETyRFsW0D9NBP = KiJFVa7Kln3PVycUSEnQNG <= l9uTQkxnOKF0VsYALlWDi; assign x1EQwZFojLp1LYxIXBaNWE = {EokQF3Q771FYsuXM046eTE, df9yw7V8ETyRFsW0D9NBP}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : y2IgBMpZH0famNY2XWfLlVH if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin upGPDbRFmGJ0jGUoSFSlo <= 5'b00000; end else begin upGPDbRFmGJ0jGUoSFSlo <= x1EQwZFojLp1LYxIXBaNWE; end end assign scXDy9YYbNjMkzYu9H6NVC = {f0Pv94BMpwnCMzWcufXc6hF, 2'b00}; assign uZFlhddYpWdV2PRdQqigiG = (df9yw7V8ETyRFsW0D9NBP == 1'b0 ? scXDy9YYbNjMkzYu9H6NVC : KiJFVa7Kln3PVycUSEnQNG); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : F1EFscGF5qvZ1uSh9OJkpG if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin SYr8j8M72olItx5mxZg3Y <= 10'b0000000000; end else begin SYr8j8M72olItx5mxZg3Y <= uZFlhddYpWdV2PRdQqigiG; end end assign ciJx9JM6wpMOOlrHHiFDNF = {SYr8j8M72olItx5mxZg3Y, 2'b01}; assign S2BiHHBn9DfCYxiINFX69C = {upGPDbRFmGJ0jGUoSFSlo, 2'b00}; assign A5VMUTy53cH6e5xVrTmqs = ({1'b0, ciJx9JM6wpMOOlrHHiFDNF}) + ({6'b0, S2BiHHBn9DfCYxiINFX69C}); assign dp2CW66DVlddH12FzsbYtB = (A5VMUTy53cH6e5xVrTmqs[12] != 1'b0 ? 12'b111111111111 : A5VMUTy53cH6e5xVrTmqs[11:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : F5Z4MbKO2IHNR1RcfbXGjH if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin LXl9oQE5X1sFOi0vAmIARG <= 32'b00000000000000000000000000000000; end else begin LXl9oQE5X1sFOi0vAmIARG <= npDxBmN6dOapdh7YCQNR6E; end end assign TaL4eG7ansmqPnA9GOrj7B = LXl9oQE5X1sFOi0vAmIARG[31:20]; assign ovy3LStQ9NhYK0h8Fs3GuF = dp2CW66DVlddH12FzsbYtB <= TaL4eG7ansmqPnA9GOrj7B; assign nFECnxinHyxo8igKFGptnB = {upGPDbRFmGJ0jGUoSFSlo, ovy3LStQ9NhYK0h8Fs3GuF}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : yRHsPlAumZ5eNVTBbdyxFG if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin QVb00VBEtaVfpEONJrgsrD <= 6'b000000; end else begin QVb00VBEtaVfpEONJrgsrD <= nFECnxinHyxo8igKFGptnB; end end assign i8Q2fmoBrZj5QeOKDTy7OXC = {SYr8j8M72olItx5mxZg3Y, 2'b00}; assign aCdbqb3Z1RZUA24wJhmb8D = (ovy3LStQ9NhYK0h8Fs3GuF == 1'b0 ? i8Q2fmoBrZj5QeOKDTy7OXC : dp2CW66DVlddH12FzsbYtB); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : hyRH3a7TEBSeUYqjyb9iuH if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin d8keq4sOv6FPsVBE0yF3SNH <= 12'b000000000000; end else begin d8keq4sOv6FPsVBE0yF3SNH <= aCdbqb3Z1RZUA24wJhmb8D; end end assign u5OcuPukOTULEzZHTQa5jE = {d8keq4sOv6FPsVBE0yF3SNH, 2'b01}; assign pnxSnkOhYHGvcrejMZZzGD = {QVb00VBEtaVfpEONJrgsrD, 2'b00}; assign pc28A478dggU3B9LCjrwKH = ({1'b0, u5OcuPukOTULEzZHTQa5jE}) + ({7'b0, pnxSnkOhYHGvcrejMZZzGD}); assign Gx4uCMMDMcZkPFg5X7j67C = (pc28A478dggU3B9LCjrwKH[14] != 1'b0 ? 14'b11111111111111 : pc28A478dggU3B9LCjrwKH[13:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : luqRHXKJ0WymWnQQiHndgC if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin VyfaXsLYCMGgAglyPOPl1C <= 32'b00000000000000000000000000000000; end else begin VyfaXsLYCMGgAglyPOPl1C <= LXl9oQE5X1sFOi0vAmIARG; end end assign Z2TjolWsiqSfSlQUx9priB = VyfaXsLYCMGgAglyPOPl1C[31:18]; assign vHqd7R6RAG8NCgLXFiRG5C = Gx4uCMMDMcZkPFg5X7j67C <= Z2TjolWsiqSfSlQUx9priB; assign j2LzkDa3ilhqsCEzuuaMJF = {QVb00VBEtaVfpEONJrgsrD, vHqd7R6RAG8NCgLXFiRG5C}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : L1bOBoyEPz6jOaW8LUHG9D if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin d8vwhmLzwzph5ZWCJmi6ErG <= 7'b0000000; end else begin d8vwhmLzwzph5ZWCJmi6ErG <= j2LzkDa3ilhqsCEzuuaMJF; end end assign POoNYqus4WpIeJLkV05T5D = {d8keq4sOv6FPsVBE0yF3SNH, 2'b00}; assign Rz1A4aD1tARfsL4hWRkGuC = (vHqd7R6RAG8NCgLXFiRG5C == 1'b0 ? POoNYqus4WpIeJLkV05T5D : Gx4uCMMDMcZkPFg5X7j67C); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : wsjaqpEBDlJnfe8pa6RvpE if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin zE0XGJgmBnFBVyzADLIUtH <= 14'b00000000000000; end else begin zE0XGJgmBnFBVyzADLIUtH <= Rz1A4aD1tARfsL4hWRkGuC; end end assign f7vtVkzvkHLoKRQDBqXTbID = {zE0XGJgmBnFBVyzADLIUtH, 2'b01}; assign xtUeqmfA0OlZnZC5um4zvE = {d8vwhmLzwzph5ZWCJmi6ErG, 2'b00}; assign l1Zuzf5TzQSJzUw3Msm6HJB = ({1'b0, f7vtVkzvkHLoKRQDBqXTbID}) + ({8'b0, xtUeqmfA0OlZnZC5um4zvE}); assign COlOv7R0Bf2iQD98SJNBZG = (l1Zuzf5TzQSJzUw3Msm6HJB[16] != 1'b0 ? 16'b1111111111111111 : l1Zuzf5TzQSJzUw3Msm6HJB[15:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : dK8Iv6LTKj9nUHsqIas7dD if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin P6kiEiTnuWYRUMrtGnBCNE <= 32'b00000000000000000000000000000000; end else begin P6kiEiTnuWYRUMrtGnBCNE <= VyfaXsLYCMGgAglyPOPl1C; end end assign xbOF64W9Ar4Lqlq1uimKrD = P6kiEiTnuWYRUMrtGnBCNE[31:16]; assign j7fDTHKDIw1b9ho08HQpp7E = COlOv7R0Bf2iQD98SJNBZG <= xbOF64W9Ar4Lqlq1uimKrD; assign as3iWC3h2hgaDUNBaZqgv = {d8vwhmLzwzph5ZWCJmi6ErG, j7fDTHKDIw1b9ho08HQpp7E}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : h88CQ12cB6YpSjrAndjy3F if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin UjnjfhzZkOwIVGTyKJXtgB <= 8'b00000000; end else begin UjnjfhzZkOwIVGTyKJXtgB <= as3iWC3h2hgaDUNBaZqgv; end end assign p5quEV42RCn3OtXuG3mHSvH = {zE0XGJgmBnFBVyzADLIUtH, 2'b00}; assign kbuD4rfjFj3gUIhRcx2cdG = (j7fDTHKDIw1b9ho08HQpp7E == 1'b0 ? p5quEV42RCn3OtXuG3mHSvH : COlOv7R0Bf2iQD98SJNBZG); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : k1CUt0kEDY8DRll3uBgCWm if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin QejN3kgI3Jo6juzY8hBlyE <= 16'b0000000000000000; end else begin QejN3kgI3Jo6juzY8hBlyE <= kbuD4rfjFj3gUIhRcx2cdG; end end assign IeHprHWybCEsl7WYUcFGsD = {QejN3kgI3Jo6juzY8hBlyE, 2'b01}; assign JIAufNDlaR5FZG2gmjhTkC = {UjnjfhzZkOwIVGTyKJXtgB, 2'b00}; assign ru0nteK8qxRvyWKiCzOgyF = ({1'b0, IeHprHWybCEsl7WYUcFGsD}) + ({9'b0, JIAufNDlaR5FZG2gmjhTkC}); assign o4ibQVfuhBHTF5NDhAQ1fKD = (ru0nteK8qxRvyWKiCzOgyF[18] != 1'b0 ? 18'b111111111111111111 : ru0nteK8qxRvyWKiCzOgyF[17:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : UBKNj7ajV0y0w8ZTet5nm if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin RtvTaElUgdpBmXzJb0yJKD <= 32'b00000000000000000000000000000000; end else begin RtvTaElUgdpBmXzJb0yJKD <= P6kiEiTnuWYRUMrtGnBCNE; end end assign MyltTFSsXFeoPojqyAjON = RtvTaElUgdpBmXzJb0yJKD[31:14]; assign hXEYb4xQxcywPjqLBUEGgD = o4ibQVfuhBHTF5NDhAQ1fKD <= MyltTFSsXFeoPojqyAjON; assign p41v0Mk0HADN0WDJBhiMxfC = {UjnjfhzZkOwIVGTyKJXtgB, hXEYb4xQxcywPjqLBUEGgD}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : kOG6Ffjkj4YAHglJQysZ6D if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin ffsa6OEyoM0DX4OPlTzw8C <= 9'b000000000; end else begin ffsa6OEyoM0DX4OPlTzw8C <= p41v0Mk0HADN0WDJBhiMxfC; end end assign nj7Uorw3TSz9rKxp2igQEC = {QejN3kgI3Jo6juzY8hBlyE, 2'b00}; assign kmD6Ilrh464BCBLVMn4VbE = (hXEYb4xQxcywPjqLBUEGgD == 1'b0 ? nj7Uorw3TSz9rKxp2igQEC : o4ibQVfuhBHTF5NDhAQ1fKD); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : B7gxnoj5znD6HTeM98beNC if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin kfbQPocRbakJ21Bwqsv0i <= 18'b000000000000000000; end else begin kfbQPocRbakJ21Bwqsv0i <= kmD6Ilrh464BCBLVMn4VbE; end end assign Iab7HeJSQoSgUz7RuhVazF = {kfbQPocRbakJ21Bwqsv0i, 2'b01}; assign jJ5plnxESkvDaAL3rZt2LB = {ffsa6OEyoM0DX4OPlTzw8C, 2'b00}; assign QEYaVcLKCNUVOqER9xXxWC = ({1'b0, Iab7HeJSQoSgUz7RuhVazF}) + ({10'b0, jJ5plnxESkvDaAL3rZt2LB}); assign pt5fnF9KyMic6eq7rU7gqD = (QEYaVcLKCNUVOqER9xXxWC[20] != 1'b0 ? 20'b11111111111111111111 : QEYaVcLKCNUVOqER9xXxWC[19:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : FVqb25uX0D3GsPefVZLTlB if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin hrT2I9W8UAX8lkCh9HwCyC <= 32'b00000000000000000000000000000000; end else begin hrT2I9W8UAX8lkCh9HwCyC <= RtvTaElUgdpBmXzJb0yJKD; end end assign cfe4isuXwwohZOaspwNnNG = hrT2I9W8UAX8lkCh9HwCyC[31:12]; assign xJZJ529nCjQslckQHtmxZH = pt5fnF9KyMic6eq7rU7gqD <= cfe4isuXwwohZOaspwNnNG; assign j7nAYb6dlFCqOFMxfcVd7QH = {ffsa6OEyoM0DX4OPlTzw8C, xJZJ529nCjQslckQHtmxZH}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : y5IVqBvXm3dThdOLiQlm2NC if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin JHUut6Rpogqw8E9skISIeG <= 10'b0000000000; end else begin JHUut6Rpogqw8E9skISIeG <= j7nAYb6dlFCqOFMxfcVd7QH; end end assign TE4W5J0afB9JODLAQ10TQF = {kfbQPocRbakJ21Bwqsv0i, 2'b00}; assign e8QGmucX9ku7ugMNMP8ZiS = (xJZJ529nCjQslckQHtmxZH == 1'b0 ? TE4W5J0afB9JODLAQ10TQF : pt5fnF9KyMic6eq7rU7gqD); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : noTZk7bnANCxfXLiopwFKB if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin gpMM7ieMx4QRfhCV7UZauE <= 20'b00000000000000000000; end else begin gpMM7ieMx4QRfhCV7UZauE <= e8QGmucX9ku7ugMNMP8ZiS; end end assign OUglDJO4thns7zNL28NuxG = {gpMM7ieMx4QRfhCV7UZauE, 2'b01}; assign C7tDtgXgfSxjvHdfE2p2hD = {JHUut6Rpogqw8E9skISIeG, 2'b00}; assign CyNDnUuxJcv2BmXf9rWncE = ({1'b0, OUglDJO4thns7zNL28NuxG}) + ({11'b0, C7tDtgXgfSxjvHdfE2p2hD}); assign MEVPG7Vi3Dy7JBBjWyUNc = (CyNDnUuxJcv2BmXf9rWncE[22] != 1'b0 ? 22'b1111111111111111111111 : CyNDnUuxJcv2BmXf9rWncE[21:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : hHqaUZt3bTf5mHLJCG9Q7 if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin azzFEVo2AvUNoNmYWBwoqH <= 32'b00000000000000000000000000000000; end else begin azzFEVo2AvUNoNmYWBwoqH <= hrT2I9W8UAX8lkCh9HwCyC; end end assign eeRMcqFduj2oNy3g1HVxSC = azzFEVo2AvUNoNmYWBwoqH[31:10]; assign jz1BZADe0coZodBEtJnz4C = MEVPG7Vi3Dy7JBBjWyUNc <= eeRMcqFduj2oNy3g1HVxSC; assign IwuuD2S9yNrHHdvvAG5YUH = {JHUut6Rpogqw8E9skISIeG, jz1BZADe0coZodBEtJnz4C}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : xijk7AdRh04whc7MH8CIGC if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin imCuL1FFwqq4jnPaCveL8E <= 11'b00000000000; end else begin imCuL1FFwqq4jnPaCveL8E <= IwuuD2S9yNrHHdvvAG5YUH; end end assign k2ck0YJnFDXHpMedhgr9qRD = {gpMM7ieMx4QRfhCV7UZauE, 2'b00}; assign sDVB7xEtvbOFj8Ui2bnoQE = (jz1BZADe0coZodBEtJnz4C == 1'b0 ? k2ck0YJnFDXHpMedhgr9qRD : MEVPG7Vi3Dy7JBBjWyUNc); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : uUsLqqhh7zC8R3Fut3SdfE if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin JVzqyten1mMc4Z5uvlfZDE <= 22'b0000000000000000000000; end else begin JVzqyten1mMc4Z5uvlfZDE <= sDVB7xEtvbOFj8Ui2bnoQE; end end assign b88drpPnD2VtwJtiEYRFQsF = {JVzqyten1mMc4Z5uvlfZDE, 2'b01}; assign qKdAaZR9hfVY5g9WEB9evF = {imCuL1FFwqq4jnPaCveL8E, 2'b00}; assign bswyonmpcfI0PoIt3aDSnF = ({1'b0, b88drpPnD2VtwJtiEYRFQsF}) + ({12'b0, qKdAaZR9hfVY5g9WEB9evF}); assign BzfSkcRvRiID6B853Sk1fE = (bswyonmpcfI0PoIt3aDSnF[24] != 1'b0 ? 24'b111111111111111111111111 : bswyonmpcfI0PoIt3aDSnF[23:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : TRt92lsaga4NyQ5SwysaxC if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin m2hoy362oakremk4ykeoJB <= 32'b00000000000000000000000000000000; end else begin m2hoy362oakremk4ykeoJB <= azzFEVo2AvUNoNmYWBwoqH; end end assign a2E5bq4xG9P8XECnOWVSMB = m2hoy362oakremk4ykeoJB[31:8]; assign s3Q2hbnFvcjqlvgMHyoBJE = BzfSkcRvRiID6B853Sk1fE <= a2E5bq4xG9P8XECnOWVSMB; assign bZEiDJSctoVjsoXa259StH = {imCuL1FFwqq4jnPaCveL8E, s3Q2hbnFvcjqlvgMHyoBJE}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : P2V9hBn0BrvUlBgRdsWO6C if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin eDBMOFTBb83n7sEEEKLXq <= 12'b000000000000; end else begin eDBMOFTBb83n7sEEEKLXq <= bZEiDJSctoVjsoXa259StH; end end assign hvkiJvP1syVDuE7eNoNFYF = {JVzqyten1mMc4Z5uvlfZDE, 2'b00}; assign cm0e9uh59eoFN2OUKptdvC = (s3Q2hbnFvcjqlvgMHyoBJE == 1'b0 ? hvkiJvP1syVDuE7eNoNFYF : BzfSkcRvRiID6B853Sk1fE); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : fV3LPZfB3qEaARITeXg9vH if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin EtkP3DOGdC8t6olD8mZndB <= 24'b000000000000000000000000; end else begin EtkP3DOGdC8t6olD8mZndB <= cm0e9uh59eoFN2OUKptdvC; end end assign iWvOu13ViXR7sawgPT1FjC = {EtkP3DOGdC8t6olD8mZndB, 2'b01}; assign FCMxV8HogSFueL98F2gNZB = {eDBMOFTBb83n7sEEEKLXq, 2'b00}; assign OqbQk3ID7Nz1GCGU2AjVl = ({1'b0, iWvOu13ViXR7sawgPT1FjC}) + ({13'b0, FCMxV8HogSFueL98F2gNZB}); assign mCdg923NHIP5asuuf0W2lH = (OqbQk3ID7Nz1GCGU2AjVl[26] != 1'b0 ? 26'b11111111111111111111111111 : OqbQk3ID7Nz1GCGU2AjVl[25:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : XetySLQTa1TDNMlT4XoQ8 if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin UWcy8pW199vG0VtRCBW2KG <= 32'b00000000000000000000000000000000; end else begin UWcy8pW199vG0VtRCBW2KG <= m2hoy362oakremk4ykeoJB; end end assign ioSpbvR6GmIfKRjNpsh2bF = UWcy8pW199vG0VtRCBW2KG[31:6]; assign WX4RpTNKBdQSVBqSWlRVFH = mCdg923NHIP5asuuf0W2lH <= ioSpbvR6GmIfKRjNpsh2bF; assign T49urcBbEEYXRINyVdZulH = {eDBMOFTBb83n7sEEEKLXq, WX4RpTNKBdQSVBqSWlRVFH}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : rjnvbHff9AyFuMs7Ecr6AC if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin e1HEl1XlshKTotIEunk6hl <= 13'b0000000000000; end else begin e1HEl1XlshKTotIEunk6hl <= T49urcBbEEYXRINyVdZulH; end end assign w7VJdxjubq01SlsqGHlxfG = {EtkP3DOGdC8t6olD8mZndB, 2'b00}; assign tTlljYwJT4O5u3alzMe2wE = (WX4RpTNKBdQSVBqSWlRVFH == 1'b0 ? w7VJdxjubq01SlsqGHlxfG : mCdg923NHIP5asuuf0W2lH); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : dBPLK3fU34jU6YX2UuU4CH if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin QPW8GtDQnJ7lqvnVJpijxF <= 26'b00000000000000000000000000; end else begin QPW8GtDQnJ7lqvnVJpijxF <= tTlljYwJT4O5u3alzMe2wE; end end assign X8nA6uSQZbaymM4A1xITNC = {QPW8GtDQnJ7lqvnVJpijxF, 2'b01}; assign iRy6kU8Izv9CM66zbzdb5E = {e1HEl1XlshKTotIEunk6hl, 2'b00}; assign KP1LyZ1AFIuavnuOnBw1VF = ({1'b0, X8nA6uSQZbaymM4A1xITNC}) + ({14'b0, iRy6kU8Izv9CM66zbzdb5E}); assign M6VKmyjZQOZXGkAKz1YjmE = (KP1LyZ1AFIuavnuOnBw1VF[28] != 1'b0 ? 28'b1111111111111111111111111111 : KP1LyZ1AFIuavnuOnBw1VF[27:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : Z9HkCRALTETLZJ6oekucLF if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin Aj7pH4hZbnjAUjVZDj9vFB <= 32'b00000000000000000000000000000000; end else begin Aj7pH4hZbnjAUjVZDj9vFB <= UWcy8pW199vG0VtRCBW2KG; end end assign DwBwYHrLgg9kBDz3J9ELdB = Aj7pH4hZbnjAUjVZDj9vFB[31:4]; assign v4mEf9URPRBLqIECbXnBDH = M6VKmyjZQOZXGkAKz1YjmE <= DwBwYHrLgg9kBDz3J9ELdB; assign NKWf6OMVvpkOpk9VSSgyRD = {e1HEl1XlshKTotIEunk6hl, v4mEf9URPRBLqIECbXnBDH}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : QogHYDEpaBJ4ySo5jnENSH if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin pQouavJJCwsKCEciQhrK3E <= 14'b00000000000000; end else begin pQouavJJCwsKCEciQhrK3E <= NKWf6OMVvpkOpk9VSSgyRD; end end assign bEAowsULkF3zy5hFKpiuSG = {QPW8GtDQnJ7lqvnVJpijxF, 2'b00}; assign yJA4o0iAYXBOPsUCeScNfC = (v4mEf9URPRBLqIECbXnBDH == 1'b0 ? bEAowsULkF3zy5hFKpiuSG : M6VKmyjZQOZXGkAKz1YjmE); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : kJvmCbdsrozdLYsfVWhN9E if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin IeN8KMSMvMg9IHSLo9n8DD <= 28'b0000000000000000000000000000; end else begin IeN8KMSMvMg9IHSLo9n8DD <= yJA4o0iAYXBOPsUCeScNfC; end end assign zJ4HWiLEv2XMiMoWf7FLPF = {IeN8KMSMvMg9IHSLo9n8DD, 2'b01}; assign AVFpT7Ib2pO9YuXeN5BZ7G = {pQouavJJCwsKCEciQhrK3E, 2'b00}; assign f7EfvG50GJ7jqsywvc9ALC = ({1'b0, zJ4HWiLEv2XMiMoWf7FLPF}) + ({15'b0, AVFpT7Ib2pO9YuXeN5BZ7G}); assign i0wZxrICRhlPz2FiwtdU8D = (f7EfvG50GJ7jqsywvc9ALC[30] != 1'b0 ? 30'b111111111111111111111111111111 : f7EfvG50GJ7jqsywvc9ALC[29:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : k9FNACRumvs3waBmRj9zhC if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin Teq2Ch748yHVvAT4uGB2FG <= 32'b00000000000000000000000000000000; end else begin Teq2Ch748yHVvAT4uGB2FG <= Aj7pH4hZbnjAUjVZDj9vFB; end end assign u5WmpPBQNytMuE3KlJIOpi = Teq2Ch748yHVvAT4uGB2FG[31:2]; assign o3K5Quha1VLfPYfrjqgd2GC = i0wZxrICRhlPz2FiwtdU8D <= u5WmpPBQNytMuE3KlJIOpi; assign i7el1SwQPx2WBbyDGEvo0HE = {pQouavJJCwsKCEciQhrK3E, o3K5Quha1VLfPYfrjqgd2GC}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : z7OkjV1u29qyU4u7w9SDePG if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin KOx599mHUoBor0KqJHxFwD <= 15'b000000000000000; end else begin KOx599mHUoBor0KqJHxFwD <= i7el1SwQPx2WBbyDGEvo0HE; end end assign faBh6P2w0PfMFOrrdKqngC = {IeN8KMSMvMg9IHSLo9n8DD, 2'b00}; assign Hh9HmtirCWU1zK1p4lc56F = (o3K5Quha1VLfPYfrjqgd2GC == 1'b0 ? faBh6P2w0PfMFOrrdKqngC : i0wZxrICRhlPz2FiwtdU8D); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : CLk3mZ7FuiHhPCS9UkW5FD if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin BqdWvf3iIjFaDgt9oYSkhG <= 30'b000000000000000000000000000000; end else begin BqdWvf3iIjFaDgt9oYSkhG <= Hh9HmtirCWU1zK1p4lc56F; end end assign SfhLiBMyxkjp1mCnRxW8FF = {BqdWvf3iIjFaDgt9oYSkhG, 2'b01}; assign BsKpUAswevf1juloThWu8D = {KOx599mHUoBor0KqJHxFwD, 2'b00}; assign RSGrktqBvyzhNztToycF6C = ({1'b0, SfhLiBMyxkjp1mCnRxW8FF}) + ({16'b0, BsKpUAswevf1juloThWu8D}); assign a3rKmat8RqcNJsLf5q2n3lF = (RSGrktqBvyzhNztToycF6C[32] != 1'b0 ? 32'b11111111111111111111111111111111 : RSGrktqBvyzhNztToycF6C[31:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : VgbxPbxi5JRL5vK69UrcMH if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin rIrurMdcINDtP7R4SI48FC <= 32'b00000000000000000000000000000000; end else begin rIrurMdcINDtP7R4SI48FC <= Teq2Ch748yHVvAT4uGB2FG; end end assign TIXiaddILO7mGZ5fWGjDCG = a3rKmat8RqcNJsLf5q2n3lF <= rIrurMdcINDtP7R4SI48FC; assign q65RX0Z30mhM7iJaeWaDrB = {KOx599mHUoBor0KqJHxFwD, TIXiaddILO7mGZ5fWGjDCG}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : Aczx50DaUmvhc1tqXErgaC if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin huOSY5XC1YM0brxFNzDqbH <= 16'b0000000000000000; end else begin huOSY5XC1YM0brxFNzDqbH <= q65RX0Z30mhM7iJaeWaDrB; end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : yqbq8XGCcWK7ainiW29o8F if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin a0r0hzxzkyJf9emryhMzNH[0] <= 16'b0000000000000000; a0r0hzxzkyJf9emryhMzNH[1] <= 16'b0000000000000000; end else begin a0r0hzxzkyJf9emryhMzNH[0] <= mSur73tREBGM65xgjFu23D[0]; a0r0hzxzkyJf9emryhMzNH[1] <= mSur73tREBGM65xgjFu23D[1]; end end assign FbFmmmgZQfWceRTyvEh1XD = a0r0hzxzkyJf9emryhMzNH[1]; assign mSur73tREBGM65xgjFu23D[0] = huOSY5XC1YM0brxFNzDqbH; assign mSur73tREBGM65xgjFu23D[1] = a0r0hzxzkyJf9emryhMzNH[0]; assign rli8whUrHAa4gMtjCDSb8G = FbFmmmgZQfWceRTyvEh1XD; assign DVmjaezJpTmh9E1RX58vDE = rli8whUrHAa4gMtjCDSb8G; assign D3zFB0T3BdpEDXphszsGdB = jQKNLtXo0Dqi6Vn3Jy2niG; assign CbG6VEOygHZYUZzB34fCPD = D3zFB0T3BdpEDXphszsGdB[31:30]; assign LRYct7GPXlUHbsVioc1vsC = 2'b01 <= CbG6VEOygHZYUZzB34fCPD; assign O5ZhenpM9MNYjlC37pcmaB = (LRYct7GPXlUHbsVioc1vsC == 1'b0 ? 1'b0 : 1'b1); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : o087uYBhztcolSYnZqD6q6C if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin VFANHQZIGPAY7b4qkN3UmC <= 1'b0; end else begin VFANHQZIGPAY7b4qkN3UmC <= O5ZhenpM9MNYjlC37pcmaB; end end assign wPuizGWKwJU15dBqzdZrBD = (LRYct7GPXlUHbsVioc1vsC == 1'b0 ? 2'b00 : 2'b01); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : jMrhiBzT6OPwwXrkyxMywG if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin mqahydaC3BSODO8RxqH5PB <= 2'b00; end else begin mqahydaC3BSODO8RxqH5PB <= wPuizGWKwJU15dBqzdZrBD; end end assign VBO1aVfkto7xu4QNiqWIZE = {mqahydaC3BSODO8RxqH5PB, 2'b01}; assign LdC0oEIcEn2u37BATOVquC = {VFANHQZIGPAY7b4qkN3UmC, 2'b00}; assign kI3sx5pDEv3shi2CwtDowE = ({1'b0, VBO1aVfkto7xu4QNiqWIZE}) + ({2'b0, LdC0oEIcEn2u37BATOVquC}); assign PHhhAthYaDH0mmviJi8guB = (kI3sx5pDEv3shi2CwtDowE[4] != 1'b0 ? 4'b1111 : kI3sx5pDEv3shi2CwtDowE[3:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : pOV9vhWMJSqNp2ULTZGgDE if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin aT9efCDUWqkTFzkLh62zcE <= 32'b00000000000000000000000000000000; end else begin aT9efCDUWqkTFzkLh62zcE <= D3zFB0T3BdpEDXphszsGdB; end end assign UNAFAbTORoRqY4QDbHcJqG = aT9efCDUWqkTFzkLh62zcE[31:28]; assign AdwV6s2RyWCMBpwC2HwLhF = PHhhAthYaDH0mmviJi8guB <= UNAFAbTORoRqY4QDbHcJqG; assign aBGGSCfHl2skiiW7NMSRqH = {VFANHQZIGPAY7b4qkN3UmC, AdwV6s2RyWCMBpwC2HwLhF}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : fg6pVoDFlEHDbvn9Bp0Vp if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin UIRrrD9huSjdHRzMx7sndE <= 2'b00; end else begin UIRrrD9huSjdHRzMx7sndE <= aBGGSCfHl2skiiW7NMSRqH; end end assign ws9KmMi5xRwv9SWSpHlEjG = {mqahydaC3BSODO8RxqH5PB, 2'b00}; assign BhAtwwns2SYFGkylFXi8BB = (AdwV6s2RyWCMBpwC2HwLhF == 1'b0 ? ws9KmMi5xRwv9SWSpHlEjG : PHhhAthYaDH0mmviJi8guB); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : r7MqoItni7FHEco0xLmTbG if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin bFIpPSFT8qi1DFuaWqyHtF <= 4'b0000; end else begin bFIpPSFT8qi1DFuaWqyHtF <= BhAtwwns2SYFGkylFXi8BB; end end assign V5pkjBsnPThxfTE1IZqGDB = {bFIpPSFT8qi1DFuaWqyHtF, 2'b01}; assign GgVTSIzPhN9ZDNsuxXlotF = {UIRrrD9huSjdHRzMx7sndE, 2'b00}; assign sPR4NMAZgx7B4yl8mD6wTF = ({1'b0, V5pkjBsnPThxfTE1IZqGDB}) + ({3'b0, GgVTSIzPhN9ZDNsuxXlotF}); assign NRJsb1CWMjRlknrudNj0vC = (sPR4NMAZgx7B4yl8mD6wTF[6] != 1'b0 ? 6'b111111 : sPR4NMAZgx7B4yl8mD6wTF[5:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : s18EYzIZosGdCVNtZ4r8NAB if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin d1GIPVaPfFgcgiwAjKvy8SG <= 32'b00000000000000000000000000000000; end else begin d1GIPVaPfFgcgiwAjKvy8SG <= aT9efCDUWqkTFzkLh62zcE; end end assign jjj0aH2qdZsn98a0jCTomE = d1GIPVaPfFgcgiwAjKvy8SG[31:26]; assign rv3m1T8mIpqw1vC5V1KXZD = NRJsb1CWMjRlknrudNj0vC <= jjj0aH2qdZsn98a0jCTomE; assign IiAS0qAOkfTGhzWxyd94bB = {UIRrrD9huSjdHRzMx7sndE, rv3m1T8mIpqw1vC5V1KXZD}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : ueOqGY2BFfy0N0E3xTecVD if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin NR1xVi9KX174l32cXe7IJE <= 3'b000; end else begin NR1xVi9KX174l32cXe7IJE <= IiAS0qAOkfTGhzWxyd94bB; end end assign lm4lGUUMg60sZsVKf4JVgB = {bFIpPSFT8qi1DFuaWqyHtF, 2'b00}; assign ivLtaKVVFqPbuQPRlcJpyD = (rv3m1T8mIpqw1vC5V1KXZD == 1'b0 ? lm4lGUUMg60sZsVKf4JVgB : NRJsb1CWMjRlknrudNj0vC); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : E23JHbq8ovefJYYVqJBZs if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin n7foXfKUGohH9shaofl43E <= 6'b000000; end else begin n7foXfKUGohH9shaofl43E <= ivLtaKVVFqPbuQPRlcJpyD; end end assign BS57yRSQtZPyqi5Bnq9psB = {n7foXfKUGohH9shaofl43E, 2'b01}; assign bJL4EEMedVetHndvDEZV5B = {NR1xVi9KX174l32cXe7IJE, 2'b00}; assign h1eiDNa2zA9F1HKjhzXOf8F = ({1'b0, BS57yRSQtZPyqi5Bnq9psB}) + ({4'b0, bJL4EEMedVetHndvDEZV5B}); assign N23SExOhay0JnnZmBL4yeF = (h1eiDNa2zA9F1HKjhzXOf8F[8] != 1'b0 ? 8'b11111111 : h1eiDNa2zA9F1HKjhzXOf8F[7:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : NWsP0VIwOBq8e43xChEK5C if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin cVgZOzpOdguVRHYqjIhuk <= 32'b00000000000000000000000000000000; end else begin cVgZOzpOdguVRHYqjIhuk <= d1GIPVaPfFgcgiwAjKvy8SG; end end assign UeTfFS2ghyunTw4P5wojCH = cVgZOzpOdguVRHYqjIhuk[31:24]; assign r2aRRQzAghfWk6CnLQvNaED = N23SExOhay0JnnZmBL4yeF <= UeTfFS2ghyunTw4P5wojCH; assign z0UZNzqu8Mq6paQqQqHK4UF = {NR1xVi9KX174l32cXe7IJE, r2aRRQzAghfWk6CnLQvNaED}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : Bp5OFRzmxd1CC496LowMeB if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin XXo1SDyBQiak88sFppTsjF <= 4'b0000; end else begin XXo1SDyBQiak88sFppTsjF <= z0UZNzqu8Mq6paQqQqHK4UF; end end assign GY9QWHEBZRjto6a1NRA3iH = {n7foXfKUGohH9shaofl43E, 2'b00}; assign zqHHk5KgIKVa1DwUKAqBXH = (r2aRRQzAghfWk6CnLQvNaED == 1'b0 ? GY9QWHEBZRjto6a1NRA3iH : N23SExOhay0JnnZmBL4yeF); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : oKKtKRNOcOmPOA82xfnvdF if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin n6lFBOQkulfdWipZ1B3mg <= 8'b00000000; end else begin n6lFBOQkulfdWipZ1B3mg <= zqHHk5KgIKVa1DwUKAqBXH; end end assign LfqJxMx8aPdx9Tg8ZpQLDE = {n6lFBOQkulfdWipZ1B3mg, 2'b01}; assign ksNnbnFsGUzsj0zxQU3sKE = {XXo1SDyBQiak88sFppTsjF, 2'b00}; assign a1iqvsOthb0rcqC3PKWRQDF = ({1'b0, LfqJxMx8aPdx9Tg8ZpQLDE}) + ({5'b0, ksNnbnFsGUzsj0zxQU3sKE}); assign YDcXhhOhmGwMKoHYiwexTC = (a1iqvsOthb0rcqC3PKWRQDF[10] != 1'b0 ? 10'b1111111111 : a1iqvsOthb0rcqC3PKWRQDF[9:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : sunv1280XLDfIINQDeYGtD if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin HA7EYu1tK22O9i8DfpQe9E <= 32'b00000000000000000000000000000000; end else begin HA7EYu1tK22O9i8DfpQe9E <= cVgZOzpOdguVRHYqjIhuk; end end assign kJiADoCkwzhBqxbx6PgBqG = HA7EYu1tK22O9i8DfpQe9E[31:22]; assign NxDv9cBGuOcye1qdzN2ZbE = YDcXhhOhmGwMKoHYiwexTC <= kJiADoCkwzhBqxbx6PgBqG; assign fkCZV6cvbAqBisxRxI0dSE = {XXo1SDyBQiak88sFppTsjF, NxDv9cBGuOcye1qdzN2ZbE}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : gGDhtGqs1i6RnFyPc1paOE if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin e0vzZybk8EaC0sU9yzfVEbH <= 5'b00000; end else begin e0vzZybk8EaC0sU9yzfVEbH <= fkCZV6cvbAqBisxRxI0dSE; end end assign KX8K4bcTmgK9iJZ4tFToED = {n6lFBOQkulfdWipZ1B3mg, 2'b00}; assign kaGb2Rgb5TMNxVjGWXMVbC = (NxDv9cBGuOcye1qdzN2ZbE == 1'b0 ? KX8K4bcTmgK9iJZ4tFToED : YDcXhhOhmGwMKoHYiwexTC); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : Mfep8NfpXDuT0AVYXpxKVB if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin c5L411ATxQWGbO5OX1TqZgH <= 10'b0000000000; end else begin c5L411ATxQWGbO5OX1TqZgH <= kaGb2Rgb5TMNxVjGWXMVbC; end end assign iR44CzvnLIWQDJIT2Bh92 = {c5L411ATxQWGbO5OX1TqZgH, 2'b01}; assign ggosYHNjNRgTTSM9nJcDSD = {e0vzZybk8EaC0sU9yzfVEbH, 2'b00}; assign z8NqtohpOQLMO57InnmOb = ({1'b0, iR44CzvnLIWQDJIT2Bh92}) + ({6'b0, ggosYHNjNRgTTSM9nJcDSD}); assign q31ojLkv58ZnYslUMTLzsC = (z8NqtohpOQLMO57InnmOb[12] != 1'b0 ? 12'b111111111111 : z8NqtohpOQLMO57InnmOb[11:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : u4VwgbZQMvzhXmEgHodv1B if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin smVaYT3RjC4ThcTM7llQyF <= 32'b00000000000000000000000000000000; end else begin smVaYT3RjC4ThcTM7llQyF <= HA7EYu1tK22O9i8DfpQe9E; end end assign p4997dIwDfgVVzHbKtpv7QF = smVaYT3RjC4ThcTM7llQyF[31:20]; assign qZOy2qjQqYVt7j2rqbDCTG = q31ojLkv58ZnYslUMTLzsC <= p4997dIwDfgVVzHbKtpv7QF; assign QoD3LztlGG71FSISslVviC = {e0vzZybk8EaC0sU9yzfVEbH, qZOy2qjQqYVt7j2rqbDCTG}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : efPXtu1Z5flWJ1wsXZezDB if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin phuPRYTWQCA8RK13saxVWH <= 6'b000000; end else begin phuPRYTWQCA8RK13saxVWH <= QoD3LztlGG71FSISslVviC; end end assign bZbQIJNhmFe85PbMpnosoE = {c5L411ATxQWGbO5OX1TqZgH, 2'b00}; assign qtXfts89aIY4wmBLUXPOB = (qZOy2qjQqYVt7j2rqbDCTG == 1'b0 ? bZbQIJNhmFe85PbMpnosoE : q31ojLkv58ZnYslUMTLzsC); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : LFOsWRAuKPhcT11o13SIIE if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin NuscntgAE20ZaRiAV7hqxC <= 12'b000000000000; end else begin NuscntgAE20ZaRiAV7hqxC <= qtXfts89aIY4wmBLUXPOB; end end assign kPLHo9hogSxDdfOl2CHNl = {NuscntgAE20ZaRiAV7hqxC, 2'b01}; assign t8xCnJCyFWgQ4D81QGbaPYD = {phuPRYTWQCA8RK13saxVWH, 2'b00}; assign pQltLIbYG2q4aRwtQURJEH = ({1'b0, kPLHo9hogSxDdfOl2CHNl}) + ({7'b0, t8xCnJCyFWgQ4D81QGbaPYD}); assign Lo0IPZ8YOZYiEHpLO42t = (pQltLIbYG2q4aRwtQURJEH[14] != 1'b0 ? 14'b11111111111111 : pQltLIbYG2q4aRwtQURJEH[13:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : jaO9zU4wDdrUEsDwH4f77D if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin x8T6JyOFCXgf5J8GjRm7OkG <= 32'b00000000000000000000000000000000; end else begin x8T6JyOFCXgf5J8GjRm7OkG <= smVaYT3RjC4ThcTM7llQyF; end end assign e9iuXqe8OquZNIsYKIaMIz = x8T6JyOFCXgf5J8GjRm7OkG[31:18]; assign HDdk8UacCG1vTeipSM5kCG = Lo0IPZ8YOZYiEHpLO42t <= e9iuXqe8OquZNIsYKIaMIz; assign B6E15sMkwvf69CPgeXdeMD = {phuPRYTWQCA8RK13saxVWH, HDdk8UacCG1vTeipSM5kCG}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : xhxyFLewOI46PjgUBkJ1BF if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin WgndoVXG1lvIDs49UGDJ6E <= 7'b0000000; end else begin WgndoVXG1lvIDs49UGDJ6E <= B6E15sMkwvf69CPgeXdeMD; end end assign pyOvyPa77c8LmSRqhL1NzC = {NuscntgAE20ZaRiAV7hqxC, 2'b00}; assign Pumm6kexkeR2FSC6LmP9s = (HDdk8UacCG1vTeipSM5kCG == 1'b0 ? pyOvyPa77c8LmSRqhL1NzC : Lo0IPZ8YOZYiEHpLO42t); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : MCHmiicPwvwEd1hLJNtGIE if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin OVKm7tgpOSGLpjnZC3LTHE <= 14'b00000000000000; end else begin OVKm7tgpOSGLpjnZC3LTHE <= Pumm6kexkeR2FSC6LmP9s; end end assign aU8NJptrwQ0dPQIyaGkVrF = {OVKm7tgpOSGLpjnZC3LTHE, 2'b01}; assign Js298tNl0lY511TfteNPUH = {WgndoVXG1lvIDs49UGDJ6E, 2'b00}; assign fQjzw0fgAbUvXvStCKuH4F = ({1'b0, aU8NJptrwQ0dPQIyaGkVrF}) + ({8'b0, Js298tNl0lY511TfteNPUH}); assign p8Ah8TzME5owYP5XfqJRi5C = (fQjzw0fgAbUvXvStCKuH4F[16] != 1'b0 ? 16'b1111111111111111 : fQjzw0fgAbUvXvStCKuH4F[15:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : GB7p60DPfnP3OP4vyMpqXG if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin w9wFocuxSkWDmPJPkThqR <= 32'b00000000000000000000000000000000; end else begin w9wFocuxSkWDmPJPkThqR <= x8T6JyOFCXgf5J8GjRm7OkG; end end assign SIrY8D5zdov6veAntRlukE = w9wFocuxSkWDmPJPkThqR[31:16]; assign DDupKb1BKahfvyZFNYIkJG = p8Ah8TzME5owYP5XfqJRi5C <= SIrY8D5zdov6veAntRlukE; assign pmpGHYek38BzarQ3qCmQrH = {WgndoVXG1lvIDs49UGDJ6E, DDupKb1BKahfvyZFNYIkJG}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : C8xIK5LDOO7EJhIuqosGl if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin JNYY5yF3xZ1TK4lLNrmXEG <= 8'b00000000; end else begin JNYY5yF3xZ1TK4lLNrmXEG <= pmpGHYek38BzarQ3qCmQrH; end end assign v7Sqzflwbh5pKJBPCHTKDEG = {OVKm7tgpOSGLpjnZC3LTHE, 2'b00}; assign IDrfZ6G75w0b2Ygh3LfQqH = (DDupKb1BKahfvyZFNYIkJG == 1'b0 ? v7Sqzflwbh5pKJBPCHTKDEG : p8Ah8TzME5owYP5XfqJRi5C); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : ial4xuqKx1PKPshVgtiNtE if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin Jddhqf0gqhZPY3wPFOoq0B <= 16'b0000000000000000; end else begin Jddhqf0gqhZPY3wPFOoq0B <= IDrfZ6G75w0b2Ygh3LfQqH; end end assign n8scxI2E0ECdA36CQrpIbcF = {Jddhqf0gqhZPY3wPFOoq0B, 2'b01}; assign d7Y8ztVAPOhsm7hvfGhOi8B = {JNYY5yF3xZ1TK4lLNrmXEG, 2'b00}; assign IowNApmWP2sledCgFHJxK = ({1'b0, n8scxI2E0ECdA36CQrpIbcF}) + ({9'b0, d7Y8ztVAPOhsm7hvfGhOi8B}); assign Sg8Rlnypyf03avWXdcL1OG = (IowNApmWP2sledCgFHJxK[18] != 1'b0 ? 18'b111111111111111111 : IowNApmWP2sledCgFHJxK[17:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : NrDYRcHyFhujXzDfa9BknE if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin XIKIDtpbTSIlhPajFWHSwG <= 32'b00000000000000000000000000000000; end else begin XIKIDtpbTSIlhPajFWHSwG <= w9wFocuxSkWDmPJPkThqR; end end assign pvJes4iUAsoX3Tn6rjCtoB = XIKIDtpbTSIlhPajFWHSwG[31:14]; assign u9XFbiauz7fSkqkXqpsNWG = Sg8Rlnypyf03avWXdcL1OG <= pvJes4iUAsoX3Tn6rjCtoB; assign w2kjxMWJYgH9lTQZFzFa1 = {JNYY5yF3xZ1TK4lLNrmXEG, u9XFbiauz7fSkqkXqpsNWG}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : Cok8kvusHMojWGnIA1nhU if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin a2rtoOfWEDzPhJ99mgT6QC <= 9'b000000000; end else begin a2rtoOfWEDzPhJ99mgT6QC <= w2kjxMWJYgH9lTQZFzFa1; end end assign wWFbZBQIqqnL6q7blY0Yb = {Jddhqf0gqhZPY3wPFOoq0B, 2'b00}; assign QIgCUQ7mCaVPNoxTkCAy2B = (u9XFbiauz7fSkqkXqpsNWG == 1'b0 ? wWFbZBQIqqnL6q7blY0Yb : Sg8Rlnypyf03avWXdcL1OG); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : NucjXndFucJOkKBEjsBkbB if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin bZ0TC5wIi5iy30a4rNIkDH <= 18'b000000000000000000; end else begin bZ0TC5wIi5iy30a4rNIkDH <= QIgCUQ7mCaVPNoxTkCAy2B; end end assign lBNV6ky8aHM84IPsYJR5n = {bZ0TC5wIi5iy30a4rNIkDH, 2'b01}; assign CncqyghSqUQTM1BqMCiVQD = {a2rtoOfWEDzPhJ99mgT6QC, 2'b00}; assign Jz4Rz7lGPIBJhH3PnjgUm = ({1'b0, lBNV6ky8aHM84IPsYJR5n}) + ({10'b0, CncqyghSqUQTM1BqMCiVQD}); assign AZ2r2El21cWt3ILZ6XvcTH = (Jz4Rz7lGPIBJhH3PnjgUm[20] != 1'b0 ? 20'b11111111111111111111 : Jz4Rz7lGPIBJhH3PnjgUm[19:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : OxraNtgTK4BUC3qX3tagYF if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin rsQbmn4FST8xbRglSdx2gB <= 32'b00000000000000000000000000000000; end else begin rsQbmn4FST8xbRglSdx2gB <= XIKIDtpbTSIlhPajFWHSwG; end end assign iDasY7iIgz0v06oml0mB = rsQbmn4FST8xbRglSdx2gB[31:12]; assign n2bWPIO8uW8vas2OgVHEQG = AZ2r2El21cWt3ILZ6XvcTH <= iDasY7iIgz0v06oml0mB; assign R6Vz9nbYsbvk5sgLGoA9gH = {a2rtoOfWEDzPhJ99mgT6QC, n2bWPIO8uW8vas2OgVHEQG}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : AQ3gquR99Sx81DcluB5H6C if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin wgs5gJPwk0LvUXsr88hTAE <= 10'b0000000000; end else begin wgs5gJPwk0LvUXsr88hTAE <= R6Vz9nbYsbvk5sgLGoA9gH; end end assign f8MC4kvmiJjXr0IW8cxs2JB = {bZ0TC5wIi5iy30a4rNIkDH, 2'b00}; assign gI1jgIcglDsIX7jWy9Max = (n2bWPIO8uW8vas2OgVHEQG == 1'b0 ? f8MC4kvmiJjXr0IW8cxs2JB : AZ2r2El21cWt3ILZ6XvcTH); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : Gwsl4835V1R3atj49yHPzC if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin qg1fRXQtNbgVxdF6yoyREF <= 20'b00000000000000000000; end else begin qg1fRXQtNbgVxdF6yoyREF <= gI1jgIcglDsIX7jWy9Max; end end assign T19dIaBYdTa9PZtZdWgMkD = {qg1fRXQtNbgVxdF6yoyREF, 2'b01}; assign GP7CX1dPzFlgdxhmIe77IC = {wgs5gJPwk0LvUXsr88hTAE, 2'b00}; assign ukHuAnhlCk8KBBDJvvXX5E = ({1'b0, T19dIaBYdTa9PZtZdWgMkD}) + ({11'b0, GP7CX1dPzFlgdxhmIe77IC}); assign WG8gzdLTcqsl8GywHjG9d = (ukHuAnhlCk8KBBDJvvXX5E[22] != 1'b0 ? 22'b1111111111111111111111 : ukHuAnhlCk8KBBDJvvXX5E[21:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : zO7cPHxbNf9FsXp6tGjAlC if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin n0NkQdqqnvMhDs423VLBKB <= 32'b00000000000000000000000000000000; end else begin n0NkQdqqnvMhDs423VLBKB <= rsQbmn4FST8xbRglSdx2gB; end end assign sTeAyrqG3sAnFH0TEwCgCC = n0NkQdqqnvMhDs423VLBKB[31:10]; assign VFMMCmH313z9JCR3kquowE = WG8gzdLTcqsl8GywHjG9d <= sTeAyrqG3sAnFH0TEwCgCC; assign z9QhOFznxLqChUzhI5cK0jG = {wgs5gJPwk0LvUXsr88hTAE, VFMMCmH313z9JCR3kquowE}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : m62Qy6fFuhoJwnTw2f3OjAD if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin DrSlN87zei4SgG4DNVrvDC <= 11'b00000000000; end else begin DrSlN87zei4SgG4DNVrvDC <= z9QhOFznxLqChUzhI5cK0jG; end end assign f7JMRjTBsPaAUm0MdIgRtnD = {qg1fRXQtNbgVxdF6yoyREF, 2'b00}; assign Xi3P8xPk5lz5vI0tMPsr6B = (VFMMCmH313z9JCR3kquowE == 1'b0 ? f7JMRjTBsPaAUm0MdIgRtnD : WG8gzdLTcqsl8GywHjG9d); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : avb95oK0VfboxLL6HWnaWB if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin f6nkTVOkasMPYCVdQ1t3RWB <= 22'b0000000000000000000000; end else begin f6nkTVOkasMPYCVdQ1t3RWB <= Xi3P8xPk5lz5vI0tMPsr6B; end end assign zjOnmfxOzwLbAed0PkfB2F = {f6nkTVOkasMPYCVdQ1t3RWB, 2'b01}; assign IfZ4i8sgfnUgsLonllpv8B = {DrSlN87zei4SgG4DNVrvDC, 2'b00}; assign E5qxoP9J21gq2LElkgURED = ({1'b0, zjOnmfxOzwLbAed0PkfB2F}) + ({12'b0, IfZ4i8sgfnUgsLonllpv8B}); assign vAlvu2utX7HZnziQ9vOxcG = (E5qxoP9J21gq2LElkgURED[24] != 1'b0 ? 24'b111111111111111111111111 : E5qxoP9J21gq2LElkgURED[23:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : N7fWNM74vwovUmLSt36rxB if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin m4y1ic6jtAcK6wabyszk2XG <= 32'b00000000000000000000000000000000; end else begin m4y1ic6jtAcK6wabyszk2XG <= n0NkQdqqnvMhDs423VLBKB; end end assign IcVjQXg4SRLKRiJxxXqZ8E = m4y1ic6jtAcK6wabyszk2XG[31:8]; assign deQ1vqISll3LmEKYH0A7SB = vAlvu2utX7HZnziQ9vOxcG <= IcVjQXg4SRLKRiJxxXqZ8E; assign c7yDah4XfUadElmPskVmLyB = {DrSlN87zei4SgG4DNVrvDC, deQ1vqISll3LmEKYH0A7SB}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : UUFsV4d6TapoO0aUdkCcwH if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin Nw9XhYz9rDGSiYWFthwTjE <= 12'b000000000000; end else begin Nw9XhYz9rDGSiYWFthwTjE <= c7yDah4XfUadElmPskVmLyB; end end assign JudNijS8FpWpflBOEYDLHG = {f6nkTVOkasMPYCVdQ1t3RWB, 2'b00}; assign b5qQKAR0z8iaZSmFCHxUOB = (deQ1vqISll3LmEKYH0A7SB == 1'b0 ? JudNijS8FpWpflBOEYDLHG : vAlvu2utX7HZnziQ9vOxcG); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : emFstOyY7NX7RAFLB7dTQD if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin jTESx94Dd1T02ZzWeEVYcF <= 24'b000000000000000000000000; end else begin jTESx94Dd1T02ZzWeEVYcF <= b5qQKAR0z8iaZSmFCHxUOB; end end assign MMf02FL20h69sCnNPkyTnG = {jTESx94Dd1T02ZzWeEVYcF, 2'b01}; assign yBpiynqDUQkwe3RYNavApF = {Nw9XhYz9rDGSiYWFthwTjE, 2'b00}; assign NOUvhKrq6oFXDc4VWYTVdC = ({1'b0, MMf02FL20h69sCnNPkyTnG}) + ({13'b0, yBpiynqDUQkwe3RYNavApF}); assign gMtX3xfic7tHemznuopkOB = (NOUvhKrq6oFXDc4VWYTVdC[26] != 1'b0 ? 26'b11111111111111111111111111 : NOUvhKrq6oFXDc4VWYTVdC[25:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : icn71kzwbSX2RlrdBCxxO if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin j4Arti1lMtcMN8FLTYwnLD <= 32'b00000000000000000000000000000000; end else begin j4Arti1lMtcMN8FLTYwnLD <= m4y1ic6jtAcK6wabyszk2XG; end end assign U2Fo3lJvtLBHW9ogfdvMME = j4Arti1lMtcMN8FLTYwnLD[31:6]; assign hTRZGt3YI59beY9UH4p1hC = gMtX3xfic7tHemznuopkOB <= U2Fo3lJvtLBHW9ogfdvMME; assign jCWS9kN2uVkHBlJLgsj6kG = {Nw9XhYz9rDGSiYWFthwTjE, hTRZGt3YI59beY9UH4p1hC}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : O0MtpKeiFYi70nmAzRwkZF if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin j02zF9SZU2kTOSADrFEpciF <= 13'b0000000000000; end else begin j02zF9SZU2kTOSADrFEpciF <= jCWS9kN2uVkHBlJLgsj6kG; end end assign c2ODxgHWlHLoVp7DmYQghEC = {jTESx94Dd1T02ZzWeEVYcF, 2'b00}; assign VZAGPjw1JyEheBnEY0qxmH = (hTRZGt3YI59beY9UH4p1hC == 1'b0 ? c2ODxgHWlHLoVp7DmYQghEC : gMtX3xfic7tHemznuopkOB); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : imrsVPCyQbyVj9j0LvqKTC if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin FEy2g40kN3tEW69WdAEGuB <= 26'b00000000000000000000000000; end else begin FEy2g40kN3tEW69WdAEGuB <= VZAGPjw1JyEheBnEY0qxmH; end end assign f7yOZ4lKvM8fXmfyUsACQD = {FEy2g40kN3tEW69WdAEGuB, 2'b01}; assign vgJ3Cr2LvuSOqY4k6A7uGE = {j02zF9SZU2kTOSADrFEpciF, 2'b00}; assign cUxMq6Y4mcjJgTtYxIGyAB = ({1'b0, f7yOZ4lKvM8fXmfyUsACQD}) + ({14'b0, vgJ3Cr2LvuSOqY4k6A7uGE}); assign xl28WnwOjU80W5ASAhe6dE = (cUxMq6Y4mcjJgTtYxIGyAB[28] != 1'b0 ? 28'b1111111111111111111111111111 : cUxMq6Y4mcjJgTtYxIGyAB[27:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : xaPB1GdeiWkBZNhQRYyBrD if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin KHqMKdR2LLNMgtSzPORlmC <= 32'b00000000000000000000000000000000; end else begin KHqMKdR2LLNMgtSzPORlmC <= j4Arti1lMtcMN8FLTYwnLD; end end assign NUD6Q6W2pS2fgKUnNEVCgD = KHqMKdR2LLNMgtSzPORlmC[31:4]; assign lg3UhZcdY7ALcP5blnn8XD = xl28WnwOjU80W5ASAhe6dE <= NUD6Q6W2pS2fgKUnNEVCgD; assign zVMIcJdSJmTolQAvSVleTE = {j02zF9SZU2kTOSADrFEpciF, lg3UhZcdY7ALcP5blnn8XD}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : L9aSEyhXHoeJgGQl0grAxH if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin kBBAFkyIMdTw9pxAjJ1PQE <= 14'b00000000000000; end else begin kBBAFkyIMdTw9pxAjJ1PQE <= zVMIcJdSJmTolQAvSVleTE; end end assign d7eCmZlCMqvmGdTJawNyWjG = {FEy2g40kN3tEW69WdAEGuB, 2'b00}; assign rIdmAf73ZEwrWcZ44F3tgH = (lg3UhZcdY7ALcP5blnn8XD == 1'b0 ? d7eCmZlCMqvmGdTJawNyWjG : xl28WnwOjU80W5ASAhe6dE); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : w8Jpzlb9Se9iys1YQQgNfE if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin bpSKi6hivc4nH6E2zzIO0F <= 28'b0000000000000000000000000000; end else begin bpSKi6hivc4nH6E2zzIO0F <= rIdmAf73ZEwrWcZ44F3tgH; end end assign jh5AUrSuZO8wqZbeaVRW2 = {bpSKi6hivc4nH6E2zzIO0F, 2'b01}; assign yhPwQJOLmQPtFG08fBKjl = {kBBAFkyIMdTw9pxAjJ1PQE, 2'b00}; assign cyg0eXE4VhRBBjgceai4dC = ({1'b0, jh5AUrSuZO8wqZbeaVRW2}) + ({15'b0, yhPwQJOLmQPtFG08fBKjl}); assign e29MWCdfscO1uEFKXjG5E = (cyg0eXE4VhRBBjgceai4dC[30] != 1'b0 ? 30'b111111111111111111111111111111 : cyg0eXE4VhRBBjgceai4dC[29:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : dF5WnZeizFpuyGR4nchPHD if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin I0k15e4Mqbps3RkfuTGQjB <= 32'b00000000000000000000000000000000; end else begin I0k15e4Mqbps3RkfuTGQjB <= KHqMKdR2LLNMgtSzPORlmC; end end assign TMGATS9eD79sBvLQD4W6iG = I0k15e4Mqbps3RkfuTGQjB[31:2]; assign WiFgj83PIvYCFc2yBQbeW = e29MWCdfscO1uEFKXjG5E <= TMGATS9eD79sBvLQD4W6iG; assign a5WzJ7XQv96wNGYwcc9tqG = {kBBAFkyIMdTw9pxAjJ1PQE, WiFgj83PIvYCFc2yBQbeW}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : VC84AGKIZTmt4vTDMtSDdF if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin ipdO2sWhLe9H5WGpausKI <= 15'b000000000000000; end else begin ipdO2sWhLe9H5WGpausKI <= a5WzJ7XQv96wNGYwcc9tqG; end end assign cIi6w7oMwXcWCEETgy8lPB = {bpSKi6hivc4nH6E2zzIO0F, 2'b00}; assign JrtSMcosjxt3HtURicDP1D = (WiFgj83PIvYCFc2yBQbeW == 1'b0 ? cIi6w7oMwXcWCEETgy8lPB : e29MWCdfscO1uEFKXjG5E); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : D2Wufo3mT6bw75XT1yjEb if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin mEmXvk5JjuKgxmWiD2PTKB <= 30'b000000000000000000000000000000; end else begin mEmXvk5JjuKgxmWiD2PTKB <= JrtSMcosjxt3HtURicDP1D; end end assign axcp60hEFY4m3CLm2qD0RF = {mEmXvk5JjuKgxmWiD2PTKB, 2'b01}; assign jkQbtWVNPA74tjUiciPhpD = {ipdO2sWhLe9H5WGpausKI, 2'b00}; assign tLOPvPysS9xFrLzWomBlzG = ({1'b0, axcp60hEFY4m3CLm2qD0RF}) + ({16'b0, jkQbtWVNPA74tjUiciPhpD}); assign v4pxjsLZ10u8ylsW5IyGeD = (tLOPvPysS9xFrLzWomBlzG[32] != 1'b0 ? 32'b11111111111111111111111111111111 : tLOPvPysS9xFrLzWomBlzG[31:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : MnQ4ILYB1z8eNnLGaLDGMC if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin AU8kfu9Bk1j6iNF7JHgrNC <= 32'b00000000000000000000000000000000; end else begin AU8kfu9Bk1j6iNF7JHgrNC <= I0k15e4Mqbps3RkfuTGQjB; end end assign adhdaT5bCy3ZoSykpu78oH = v4pxjsLZ10u8ylsW5IyGeD <= AU8kfu9Bk1j6iNF7JHgrNC; assign kmeXG1ZdV7nLMdzktaC88C = {ipdO2sWhLe9H5WGpausKI, adhdaT5bCy3ZoSykpu78oH}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : Ue5dCY18D5c90IhdvwRlvB if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin oBIxcPTGR95iZNFbr4227G <= 16'b0000000000000000; end else begin oBIxcPTGR95iZNFbr4227G <= kmeXG1ZdV7nLMdzktaC88C; end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : qrGDgS8OUwXdApQx8AuPeF if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin s16lp7vAtcFZ2wwPaIkgzB[0] <= 16'b0000000000000000; s16lp7vAtcFZ2wwPaIkgzB[1] <= 16'b0000000000000000; end else begin s16lp7vAtcFZ2wwPaIkgzB[0] <= QH69kVWWgj2WJadmvpUaPF[0]; s16lp7vAtcFZ2wwPaIkgzB[1] <= QH69kVWWgj2WJadmvpUaPF[1]; end end assign FS8ak02sQNsotNaSejJzOF = s16lp7vAtcFZ2wwPaIkgzB[1]; assign QH69kVWWgj2WJadmvpUaPF[0] = oBIxcPTGR95iZNFbr4227G; assign QH69kVWWgj2WJadmvpUaPF[1] = s16lp7vAtcFZ2wwPaIkgzB[0]; assign s7iMbfZ00UZszqLEi06wYE = FS8ak02sQNsotNaSejJzOF; assign c50jzfprXP85SKSfjge64NC = s7iMbfZ00UZszqLEi06wYE; assign YAPbE5XIglo6YQglskaaWD = rosLsgtHKD6hJ64eM2pegF; assign b4c80DCXt5syU5YZsPFg8fG = YAPbE5XIglo6YQglskaaWD[31:30]; assign aeA4SROkYBwZ6Vg6wePll = 2'b01 <= b4c80DCXt5syU5YZsPFg8fG; assign VLU8KlCAVdk3z1akf8lgXG = (aeA4SROkYBwZ6Vg6wePll == 1'b0 ? 1'b0 : 1'b1); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : zmlqh5ak7QvPAi5I1knNwE if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin b00qa2rJFIB1ZMqONGFopXG <= 1'b0; end else begin b00qa2rJFIB1ZMqONGFopXG <= VLU8KlCAVdk3z1akf8lgXG; end end assign xmRFmcImcIZ7hAGSB5Bu8E = (aeA4SROkYBwZ6Vg6wePll == 1'b0 ? 2'b00 : 2'b01); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : OC0Y23ntcq84h1w0tW31o if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin SKbN7GhZfEspFZRKIkIVmF <= 2'b00; end else begin SKbN7GhZfEspFZRKIkIVmF <= xmRFmcImcIZ7hAGSB5Bu8E; end end assign Js5jS7mG04lv6SG081bBdD = {SKbN7GhZfEspFZRKIkIVmF, 2'b01}; assign n1zMPjaeIWPwBCg7gfpFRw = {b00qa2rJFIB1ZMqONGFopXG, 2'b00}; assign JSVnqT7wQsMpSEZncqnKU = ({1'b0, Js5jS7mG04lv6SG081bBdD}) + ({2'b0, n1zMPjaeIWPwBCg7gfpFRw}); assign d8YQiHX7vIPrjtzcNsFfqUC = (JSVnqT7wQsMpSEZncqnKU[4] != 1'b0 ? 4'b1111 : JSVnqT7wQsMpSEZncqnKU[3:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : js2usPMTsyWpKovYxVezTG if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin PkXpzwBbQLQYvzhTqlk7wB <= 32'b00000000000000000000000000000000; end else begin PkXpzwBbQLQYvzhTqlk7wB <= YAPbE5XIglo6YQglskaaWD; end end assign w7Sh4wi1uZ8tdPQjGm2IyBB = PkXpzwBbQLQYvzhTqlk7wB[31:28]; assign JIk51ZYgI4bjmkaz1s3ocD = d8YQiHX7vIPrjtzcNsFfqUC <= w7Sh4wi1uZ8tdPQjGm2IyBB; assign p5vFo8g1m0abgHiHdIbMIB = {b00qa2rJFIB1ZMqONGFopXG, JIk51ZYgI4bjmkaz1s3ocD}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : HbtXBgraohek4ykc27jTLH if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin nNsb6XV1QdVOT8po6E0QRC <= 2'b00; end else begin nNsb6XV1QdVOT8po6E0QRC <= p5vFo8g1m0abgHiHdIbMIB; end end assign f2eRR8CFkJiACbGc7JLrHC = {SKbN7GhZfEspFZRKIkIVmF, 2'b00}; assign m2es1PMsJ2xQuYLiPnHr1 = (JIk51ZYgI4bjmkaz1s3ocD == 1'b0 ? f2eRR8CFkJiACbGc7JLrHC : d8YQiHX7vIPrjtzcNsFfqUC); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : iSFI4s6KUprLOPZMXEA6sC if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin UGlnA3qCFkn9R10JNKEmWB <= 4'b0000; end else begin UGlnA3qCFkn9R10JNKEmWB <= m2es1PMsJ2xQuYLiPnHr1; end end assign f7i6sgURXoacv9zlCx7k8pE = {UGlnA3qCFkn9R10JNKEmWB, 2'b01}; assign gFnPRfLYr5mEttAuZT5TNG = {nNsb6XV1QdVOT8po6E0QRC, 2'b00}; assign AFbX6YpTqq1eBEyQFqseMC = ({1'b0, f7i6sgURXoacv9zlCx7k8pE}) + ({3'b0, gFnPRfLYr5mEttAuZT5TNG}); assign qqZdHvncdEpi1f3UX3FiLH = (AFbX6YpTqq1eBEyQFqseMC[6] != 1'b0 ? 6'b111111 : AFbX6YpTqq1eBEyQFqseMC[5:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : RxteYmlEqdldcuNsOtYO5F if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin Pz7nVzONTu3jrA61HPdb5G <= 32'b00000000000000000000000000000000; end else begin Pz7nVzONTu3jrA61HPdb5G <= PkXpzwBbQLQYvzhTqlk7wB; end end assign cr5TMAj7bawp4OzGhelvYC = Pz7nVzONTu3jrA61HPdb5G[31:26]; assign uSBJDL0TF4CJ5LqsokDLtC = qqZdHvncdEpi1f3UX3FiLH <= cr5TMAj7bawp4OzGhelvYC; assign FDrOrbrGZpLR2snFBNYfgG = {nNsb6XV1QdVOT8po6E0QRC, uSBJDL0TF4CJ5LqsokDLtC}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : J406hUZKHTolEnc8TL4A2G if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin y1AuRFIyn548BXgwQF0sZdE <= 3'b000; end else begin y1AuRFIyn548BXgwQF0sZdE <= FDrOrbrGZpLR2snFBNYfgG; end end assign U6ZX5GALoV26phzqBZLxwB = {UGlnA3qCFkn9R10JNKEmWB, 2'b00}; assign lEpIUGd5Cr0vd5frOPY3ZB = (uSBJDL0TF4CJ5LqsokDLtC == 1'b0 ? U6ZX5GALoV26phzqBZLxwB : qqZdHvncdEpi1f3UX3FiLH); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : c7sKzB5s7u26W2Twm2181F if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin Y1kJ6m5YlbS5HZjCnkaC1D <= 6'b000000; end else begin Y1kJ6m5YlbS5HZjCnkaC1D <= lEpIUGd5Cr0vd5frOPY3ZB; end end assign OsCJQX96BJolsZ5d0oBzoG = {Y1kJ6m5YlbS5HZjCnkaC1D, 2'b01}; assign MXb346opbIN11K8xrTYv0F = {y1AuRFIyn548BXgwQF0sZdE, 2'b00}; assign JiuDBTKkk3DmNTKhQeVyEE = ({1'b0, OsCJQX96BJolsZ5d0oBzoG}) + ({4'b0, MXb346opbIN11K8xrTYv0F}); assign cepH0TZ1Fi8TpQGwHx2WYE = (JiuDBTKkk3DmNTKhQeVyEE[8] != 1'b0 ? 8'b11111111 : JiuDBTKkk3DmNTKhQeVyEE[7:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : nIIolWZus0eZh1pRW6q2QG if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin cUOLCqZop1yocpR9PH5jiF <= 32'b00000000000000000000000000000000; end else begin cUOLCqZop1yocpR9PH5jiF <= Pz7nVzONTu3jrA61HPdb5G; end end assign Y8QYTUsOLW2ORrnUf75Vg = cUOLCqZop1yocpR9PH5jiF[31:24]; assign mRBRsCt0Pgu3ZY8PRCi0oD = cepH0TZ1Fi8TpQGwHx2WYE <= Y8QYTUsOLW2ORrnUf75Vg; assign n4tG0JS2MvMz1aVTykyRDpD = {y1AuRFIyn548BXgwQF0sZdE, mRBRsCt0Pgu3ZY8PRCi0oD}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : jomD4t3KmJ0iN3CWDkV0kC if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin CI6B2HVMFRzDx37oEWjIuE <= 4'b0000; end else begin CI6B2HVMFRzDx37oEWjIuE <= n4tG0JS2MvMz1aVTykyRDpD; end end assign VSMVYe1a2T37zL1SHKrC2G = {Y1kJ6m5YlbS5HZjCnkaC1D, 2'b00}; assign w2M0mYanih9pVwcHbeGmhkC = (mRBRsCt0Pgu3ZY8PRCi0oD == 1'b0 ? VSMVYe1a2T37zL1SHKrC2G : cepH0TZ1Fi8TpQGwHx2WYE); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : pecE1fGeY9jBzvW60omnnC if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin x08SSTqzuST0npo22yvHD1 <= 8'b00000000; end else begin x08SSTqzuST0npo22yvHD1 <= w2M0mYanih9pVwcHbeGmhkC; end end assign NrGTCqt9rkin8JxxJzivMC = {x08SSTqzuST0npo22yvHD1, 2'b01}; assign sMUm3XDWkY9euUemzzSHsD = {CI6B2HVMFRzDx37oEWjIuE, 2'b00}; assign qjrpTJyWev1g925QNDAW1F = ({1'b0, NrGTCqt9rkin8JxxJzivMC}) + ({5'b0, sMUm3XDWkY9euUemzzSHsD}); assign SFmRqM1SKlq0XxdjenL8yC = (qjrpTJyWev1g925QNDAW1F[10] != 1'b0 ? 10'b1111111111 : qjrpTJyWev1g925QNDAW1F[9:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : i2F6fouwQT1llaBiDx1IKyE if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin darCJM0vPSpQ6IgQNZHgPC <= 32'b00000000000000000000000000000000; end else begin darCJM0vPSpQ6IgQNZHgPC <= cUOLCqZop1yocpR9PH5jiF; end end assign YQ3g2H8nF3dqmEyVDvXGRD = darCJM0vPSpQ6IgQNZHgPC[31:22]; assign PSPwNHQ13FhdLM6OMJRHmB = SFmRqM1SKlq0XxdjenL8yC <= YQ3g2H8nF3dqmEyVDvXGRD; assign NQ4pAf9vZ8Xx4lGiiOXU6D = {CI6B2HVMFRzDx37oEWjIuE, PSPwNHQ13FhdLM6OMJRHmB}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : HwFAZ1JsOb41uOOEH8lkcE if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin sJ6GWhkNdag4yzDVnIXRZE <= 5'b00000; end else begin sJ6GWhkNdag4yzDVnIXRZE <= NQ4pAf9vZ8Xx4lGiiOXU6D; end end assign ObGqdHNTbg4VcYpEbgQjKB = {x08SSTqzuST0npo22yvHD1, 2'b00}; assign DRHq6AFeMUbFXJu9ozWhfD = (PSPwNHQ13FhdLM6OMJRHmB == 1'b0 ? ObGqdHNTbg4VcYpEbgQjKB : SFmRqM1SKlq0XxdjenL8yC); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : LFdRYQD7d8GtK76HWDkXSB if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin aAlJVECF2UJ0il926uH1xF <= 10'b0000000000; end else begin aAlJVECF2UJ0il926uH1xF <= DRHq6AFeMUbFXJu9ozWhfD; end end assign y1txMzBbEmvxmMKJpM7J1iB = {aAlJVECF2UJ0il926uH1xF, 2'b01}; assign wSKM2kCYmT1b8JpcHR77rE = {sJ6GWhkNdag4yzDVnIXRZE, 2'b00}; assign p3FlB7G5wQcEKEanZhV9aF = ({1'b0, y1txMzBbEmvxmMKJpM7J1iB}) + ({6'b0, wSKM2kCYmT1b8JpcHR77rE}); assign v4aA671Zjc8PT2J1KV8nzkD = (p3FlB7G5wQcEKEanZhV9aF[12] != 1'b0 ? 12'b111111111111 : p3FlB7G5wQcEKEanZhV9aF[11:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : LFLQSkFglj6R7HRnaAXTI if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin URZZIGLG4aIgBvyK6bwvuF <= 32'b00000000000000000000000000000000; end else begin URZZIGLG4aIgBvyK6bwvuF <= darCJM0vPSpQ6IgQNZHgPC; end end assign q92Pz7xfru0n25cOdhefGB = URZZIGLG4aIgBvyK6bwvuF[31:20]; assign nqCCuMllPTQCxAwb4BAHtF = v4aA671Zjc8PT2J1KV8nzkD <= q92Pz7xfru0n25cOdhefGB; assign m2Xf3fQbkf2EKah6ia1rhrB = {sJ6GWhkNdag4yzDVnIXRZE, nqCCuMllPTQCxAwb4BAHtF}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : ptiPOPo4VRWr8xDjmSaKQB if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin DP1rxfHwjNcmCS5dP7UEvH <= 6'b000000; end else begin DP1rxfHwjNcmCS5dP7UEvH <= m2Xf3fQbkf2EKah6ia1rhrB; end end assign In2u3aBla1oHkNHMApLKsH = {aAlJVECF2UJ0il926uH1xF, 2'b00}; assign RhvWLtfm9kbIPah6Xmhz5B = (nqCCuMllPTQCxAwb4BAHtF == 1'b0 ? In2u3aBla1oHkNHMApLKsH : v4aA671Zjc8PT2J1KV8nzkD); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : k7PJBBs55VLk9SWwhJGAaUH if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin ulxawSs2t7mfLDUIwzjgMH <= 12'b000000000000; end else begin ulxawSs2t7mfLDUIwzjgMH <= RhvWLtfm9kbIPah6Xmhz5B; end end assign QogFm8TTkYvdd1pOETS8GE = {ulxawSs2t7mfLDUIwzjgMH, 2'b01}; assign odys5fwKXDkTPl2xGW5md = {DP1rxfHwjNcmCS5dP7UEvH, 2'b00}; assign jUoV3u5hOQ3V3P9X4L422G = ({1'b0, QogFm8TTkYvdd1pOETS8GE}) + ({7'b0, odys5fwKXDkTPl2xGW5md}); assign lKy8gFEyss6k09Lab0TIyD = (jUoV3u5hOQ3V3P9X4L422G[14] != 1'b0 ? 14'b11111111111111 : jUoV3u5hOQ3V3P9X4L422G[13:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : MOqMsQk0UftMXTXxLbDEmF if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin o9IXOBjy3eJadOxzwMZYCD <= 32'b00000000000000000000000000000000; end else begin o9IXOBjy3eJadOxzwMZYCD <= URZZIGLG4aIgBvyK6bwvuF; end end assign afhwDwKsffj7ws30MIdif = o9IXOBjy3eJadOxzwMZYCD[31:18]; assign gzAMKqGsdPMTGqF8e9aodB = lKy8gFEyss6k09Lab0TIyD <= afhwDwKsffj7ws30MIdif; assign vMT5nzjGBRaywF0w7bpHnH = {DP1rxfHwjNcmCS5dP7UEvH, gzAMKqGsdPMTGqF8e9aodB}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : cDFjfvlUF0fZKMdf3bhVM if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin kQOxLlINqlKIXn0R43wTvH <= 7'b0000000; end else begin kQOxLlINqlKIXn0R43wTvH <= vMT5nzjGBRaywF0w7bpHnH; end end assign GIyfilklKRkkteItBi4jVG = {ulxawSs2t7mfLDUIwzjgMH, 2'b00}; assign cDG7Ga2x2ulXJ9HZ0kU6XE = (gzAMKqGsdPMTGqF8e9aodB == 1'b0 ? GIyfilklKRkkteItBi4jVG : lKy8gFEyss6k09Lab0TIyD); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : lhpHHWirIwICfpenrkCiLC if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin cOQeVrl2Kc2AaEV3A3SKVB <= 14'b00000000000000; end else begin cOQeVrl2Kc2AaEV3A3SKVB <= cDG7Ga2x2ulXJ9HZ0kU6XE; end end assign oUr9Z0wSJ8NEbpWbUr40O = {cOQeVrl2Kc2AaEV3A3SKVB, 2'b01}; assign v99YLq8JtK6czSdvv7sUwZH = {kQOxLlINqlKIXn0R43wTvH, 2'b00}; assign OlUTROE94KsCPuYIZdRVnD = ({1'b0, oUr9Z0wSJ8NEbpWbUr40O}) + ({8'b0, v99YLq8JtK6czSdvv7sUwZH}); assign q2d5CtZFCBdgowZqGzc7c = (OlUTROE94KsCPuYIZdRVnD[16] != 1'b0 ? 16'b1111111111111111 : OlUTROE94KsCPuYIZdRVnD[15:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : ZfSYbwyt4lND1qQcN7ycbE if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin XMliVuWBVwOcOPEdVe2sbD <= 32'b00000000000000000000000000000000; end else begin XMliVuWBVwOcOPEdVe2sbD <= o9IXOBjy3eJadOxzwMZYCD; end end assign H7HCojLu6xl0FDsspFgeF = XMliVuWBVwOcOPEdVe2sbD[31:16]; assign V5HChjE9NVsTIubsNiixTD = q2d5CtZFCBdgowZqGzc7c <= H7HCojLu6xl0FDsspFgeF; assign r0fdrd8QpMOua7OUDgRkvlE = {kQOxLlINqlKIXn0R43wTvH, V5HChjE9NVsTIubsNiixTD}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : gJUIP3z3HTn2lwFeHamzBF if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin ziHkTpSLxytlkstnKqPgtD <= 8'b00000000; end else begin ziHkTpSLxytlkstnKqPgtD <= r0fdrd8QpMOua7OUDgRkvlE; end end assign TrSsPsucRJCHZyiwqiAxYG = {cOQeVrl2Kc2AaEV3A3SKVB, 2'b00}; assign Bbz9EGUOWN194RSqeY9vzE = (V5HChjE9NVsTIubsNiixTD == 1'b0 ? TrSsPsucRJCHZyiwqiAxYG : q2d5CtZFCBdgowZqGzc7c); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : C8wgiHAOChFamV2RfbSbE if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin P41QmEa2IVlG6Gw1uNCuYC <= 16'b0000000000000000; end else begin P41QmEa2IVlG6Gw1uNCuYC <= Bbz9EGUOWN194RSqeY9vzE; end end assign liAyj9i3OaG5qj3ww4zBjB = {P41QmEa2IVlG6Gw1uNCuYC, 2'b01}; assign yCyP1ziVlDiJpYzdd6YPVG = {ziHkTpSLxytlkstnKqPgtD, 2'b00}; assign arTIxO8ttVfgZOyW4PzlzC = ({1'b0, liAyj9i3OaG5qj3ww4zBjB}) + ({9'b0, yCyP1ziVlDiJpYzdd6YPVG}); assign dCaoI2qtg6pmjm3MVxzJKH = (arTIxO8ttVfgZOyW4PzlzC[18] != 1'b0 ? 18'b111111111111111111 : arTIxO8ttVfgZOyW4PzlzC[17:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : G0iL9dsuBZff3W5VETWJmB if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin dCOpIGH8phIdHUSJlDSfvG <= 32'b00000000000000000000000000000000; end else begin dCOpIGH8phIdHUSJlDSfvG <= XMliVuWBVwOcOPEdVe2sbD; end end assign oflUhi5A8v1YWG7yE5g8i = dCOpIGH8phIdHUSJlDSfvG[31:14]; assign g93FJ0IBN4c66etyHmEs3zG = dCaoI2qtg6pmjm3MVxzJKH <= oflUhi5A8v1YWG7yE5g8i; assign OeVgNvqOmoHvuonJYQ60DE = {ziHkTpSLxytlkstnKqPgtD, g93FJ0IBN4c66etyHmEs3zG}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : FibD9MbfNFrMguvmD6KpHG if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin zQDpOsty76yxOjWPsK2jX <= 9'b000000000; end else begin zQDpOsty76yxOjWPsK2jX <= OeVgNvqOmoHvuonJYQ60DE; end end assign OnMuHOtaSmv6vr0BtqpDUB = {P41QmEa2IVlG6Gw1uNCuYC, 2'b00}; assign h3EKSUN8gsftz7jQO1rdxBE = (g93FJ0IBN4c66etyHmEs3zG == 1'b0 ? OnMuHOtaSmv6vr0BtqpDUB : dCaoI2qtg6pmjm3MVxzJKH); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : ykZUeIdLsFE36blN5bFJYH if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin Dgv0nOPwuFJGc4GAqTimbH <= 18'b000000000000000000; end else begin Dgv0nOPwuFJGc4GAqTimbH <= h3EKSUN8gsftz7jQO1rdxBE; end end assign woO6WUPEUZHhCxslCmpXsD = {Dgv0nOPwuFJGc4GAqTimbH, 2'b01}; assign n6flnvH1JRdcq5tHRAY4lC = {zQDpOsty76yxOjWPsK2jX, 2'b00}; assign Y4ORnDxB7EutyM3R3AYoLF = ({1'b0, woO6WUPEUZHhCxslCmpXsD}) + ({10'b0, n6flnvH1JRdcq5tHRAY4lC}); assign kpoCQdFe8llOB4VroSkRWB = (Y4ORnDxB7EutyM3R3AYoLF[20] != 1'b0 ? 20'b11111111111111111111 : Y4ORnDxB7EutyM3R3AYoLF[19:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : eaNeGxELd8oN8Uk74x9RwF if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin WpoaYGV1NzHQJMT5jm5HyC <= 32'b00000000000000000000000000000000; end else begin WpoaYGV1NzHQJMT5jm5HyC <= dCOpIGH8phIdHUSJlDSfvG; end end assign p5ZR7b2BqOcgrhqd260UTF = WpoaYGV1NzHQJMT5jm5HyC[31:12]; assign G44bIdnYp2VbJFdrHB9ZC = kpoCQdFe8llOB4VroSkRWB <= p5ZR7b2BqOcgrhqd260UTF; assign ZWAF6ra3GkzT56Oefe3NLF = {zQDpOsty76yxOjWPsK2jX, G44bIdnYp2VbJFdrHB9ZC}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : yQQRjFHHzq9QffBstTuUzC if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin ATgyH1zIQ4sJ6Hz7GqMsCF <= 10'b0000000000; end else begin ATgyH1zIQ4sJ6Hz7GqMsCF <= ZWAF6ra3GkzT56Oefe3NLF; end end assign lIdXhiWJIC9ldEsDa0NXZE = {Dgv0nOPwuFJGc4GAqTimbH, 2'b00}; assign P90P58Xa7n44tjlKivSZ8 = (G44bIdnYp2VbJFdrHB9ZC == 1'b0 ? lIdXhiWJIC9ldEsDa0NXZE : kpoCQdFe8llOB4VroSkRWB); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : WjebgxbXfkFId7gqZkwzuB if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin gyufbtlPcbpsc3XTEswKdB <= 20'b00000000000000000000; end else begin gyufbtlPcbpsc3XTEswKdB <= P90P58Xa7n44tjlKivSZ8; end end assign H7hJJQFtPQpIus6wdn7lu = {gyufbtlPcbpsc3XTEswKdB, 2'b01}; assign jCUl3tPIcmmqDiSckg2hhD = {ATgyH1zIQ4sJ6Hz7GqMsCF, 2'b00}; assign wIaIyn7lrKf0kblWE9XkjC = ({1'b0, H7hJJQFtPQpIus6wdn7lu}) + ({11'b0, jCUl3tPIcmmqDiSckg2hhD}); assign fFumSIcnLnWln2qYLinPuE = (wIaIyn7lrKf0kblWE9XkjC[22] != 1'b0 ? 22'b1111111111111111111111 : wIaIyn7lrKf0kblWE9XkjC[21:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : nU3uqZPVV7BZYGEQgW51a if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin nRdqcvDbm319JQcsXwul4F <= 32'b00000000000000000000000000000000; end else begin nRdqcvDbm319JQcsXwul4F <= WpoaYGV1NzHQJMT5jm5HyC; end end assign m7vHNxrFnoDjp1IrlzZ9fQB = nRdqcvDbm319JQcsXwul4F[31:10]; assign QYXTpn7JNO59MwFJCQmpxG = fFumSIcnLnWln2qYLinPuE <= m7vHNxrFnoDjp1IrlzZ9fQB; assign Dx1qecvaNRk0C8Sp1BRC7E = {ATgyH1zIQ4sJ6Hz7GqMsCF, QYXTpn7JNO59MwFJCQmpxG}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : XgNUiGOXNFpgFTVjMNUgvG if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin YJM4uTYV0GNEIq6Ts1WqdG <= 11'b00000000000; end else begin YJM4uTYV0GNEIq6Ts1WqdG <= Dx1qecvaNRk0C8Sp1BRC7E; end end assign u8NrYi3OMqbhK9yByGZs9PB = {gyufbtlPcbpsc3XTEswKdB, 2'b00}; assign rwO0PhKT8dAkniV0s365fH = (QYXTpn7JNO59MwFJCQmpxG == 1'b0 ? u8NrYi3OMqbhK9yByGZs9PB : fFumSIcnLnWln2qYLinPuE); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : RfQvgqALibFxy3FFlFqEb if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin QEFCsmo4y0LLYuDoykR98B <= 22'b0000000000000000000000; end else begin QEFCsmo4y0LLYuDoykR98B <= rwO0PhKT8dAkniV0s365fH; end end assign RX0sHsM1Nzw8rn3ouqfTE = {QEFCsmo4y0LLYuDoykR98B, 2'b01}; assign uiKvXhWqzaIyVELDYBl2pC = {YJM4uTYV0GNEIq6Ts1WqdG, 2'b00}; assign VpP6fnKzcKN32HJtlCGIuD = ({1'b0, RX0sHsM1Nzw8rn3ouqfTE}) + ({12'b0, uiKvXhWqzaIyVELDYBl2pC}); assign e3PfhueHdzlIuEVJBllUSi = (VpP6fnKzcKN32HJtlCGIuD[24] != 1'b0 ? 24'b111111111111111111111111 : VpP6fnKzcKN32HJtlCGIuD[23:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : guoYmWVLvRTjtWv6EHUXAF if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin PQtoGuipN4OobbDKTpW4zB <= 32'b00000000000000000000000000000000; end else begin PQtoGuipN4OobbDKTpW4zB <= nRdqcvDbm319JQcsXwul4F; end end assign kvSoFz62JUu4jx44u4ZCsC = PQtoGuipN4OobbDKTpW4zB[31:8]; assign vg0CbYzueQThdby6EnMwrC = e3PfhueHdzlIuEVJBllUSi <= kvSoFz62JUu4jx44u4ZCsC; assign gCzr56bCiioiPJ7vxpKGRE = {YJM4uTYV0GNEIq6Ts1WqdG, vg0CbYzueQThdby6EnMwrC}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : Z5eCAKHpl8XtSqvEHMNdlB if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin g1i4ElfCXQ9sMqQ8agpYlLC <= 12'b000000000000; end else begin g1i4ElfCXQ9sMqQ8agpYlLC <= gCzr56bCiioiPJ7vxpKGRE; end end assign TrlkOR4z072dMOyjD8yJtE = {QEFCsmo4y0LLYuDoykR98B, 2'b00}; assign pDEdPRJUIcsUQQ8UmXGdJH = (vg0CbYzueQThdby6EnMwrC == 1'b0 ? TrlkOR4z072dMOyjD8yJtE : e3PfhueHdzlIuEVJBllUSi); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : JSLDzXj40Ko2lf4IYQWfCH if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin s85203G8LCtqp2Q4Hln8eDD <= 24'b000000000000000000000000; end else begin s85203G8LCtqp2Q4Hln8eDD <= pDEdPRJUIcsUQQ8UmXGdJH; end end assign voKrZH4np5NWTctmsz4oFH = {s85203G8LCtqp2Q4Hln8eDD, 2'b01}; assign e1Rl7kcQNObhKfOXtWutrG = {g1i4ElfCXQ9sMqQ8agpYlLC, 2'b00}; assign Taj7HNFKppS43yrU3qKE1B = ({1'b0, voKrZH4np5NWTctmsz4oFH}) + ({13'b0, e1Rl7kcQNObhKfOXtWutrG}); assign L3nPxZVh5u3VVA1rdbb4QC = (Taj7HNFKppS43yrU3qKE1B[26] != 1'b0 ? 26'b11111111111111111111111111 : Taj7HNFKppS43yrU3qKE1B[25:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : i2I5hfPC0jXxTg8KfEPfOaC if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin DqFCXgxzTWTDDQbslRF6E <= 32'b00000000000000000000000000000000; end else begin DqFCXgxzTWTDDQbslRF6E <= PQtoGuipN4OobbDKTpW4zB; end end assign d3KDtpVH3H0bcfiybpzeSnB = DqFCXgxzTWTDDQbslRF6E[31:6]; assign sGiOEpItJbE2kz8n13WEwF = L3nPxZVh5u3VVA1rdbb4QC <= d3KDtpVH3H0bcfiybpzeSnB; assign zFwPpMKHPaoWNlMcn3Ooz = {g1i4ElfCXQ9sMqQ8agpYlLC, sGiOEpItJbE2kz8n13WEwF}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : LOXkliCZx7hktP0H2as1SB if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin L8G5zN2h3nNrCok5TCsJbE <= 13'b0000000000000; end else begin L8G5zN2h3nNrCok5TCsJbE <= zFwPpMKHPaoWNlMcn3Ooz; end end assign BOaYPwGg4vIF3dmZHl7rWE = {s85203G8LCtqp2Q4Hln8eDD, 2'b00}; assign IJwTxkeWtn7iKzAUHVUPeH = (sGiOEpItJbE2kz8n13WEwF == 1'b0 ? BOaYPwGg4vIF3dmZHl7rWE : L3nPxZVh5u3VVA1rdbb4QC); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : JAPfvQyedaFSPQAoARrAQB if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin DXqu7TpZsKBJkGAUCIfEdB <= 26'b00000000000000000000000000; end else begin DXqu7TpZsKBJkGAUCIfEdB <= IJwTxkeWtn7iKzAUHVUPeH; end end assign wxD3MMuIUYxbh5lNx5wYZE = {DXqu7TpZsKBJkGAUCIfEdB, 2'b01}; assign sIVqloL9MjkDXMyZqNgFi = {L8G5zN2h3nNrCok5TCsJbE, 2'b00}; assign R5FT4wZn7DjE5FtgHFUm3E = ({1'b0, wxD3MMuIUYxbh5lNx5wYZE}) + ({14'b0, sIVqloL9MjkDXMyZqNgFi}); assign on0J0v1C0T4Vx5BAyNciCG = (R5FT4wZn7DjE5FtgHFUm3E[28] != 1'b0 ? 28'b1111111111111111111111111111 : R5FT4wZn7DjE5FtgHFUm3E[27:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : nX3kjnvIKGzATz9y6uXbKF if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin zjMYjjAxK45sdDEQ0XFXOG <= 32'b00000000000000000000000000000000; end else begin zjMYjjAxK45sdDEQ0XFXOG <= DqFCXgxzTWTDDQbslRF6E; end end assign xbDZHFjT9czSWoXqDrDalH = zjMYjjAxK45sdDEQ0XFXOG[31:4]; assign rIIATJviRgNIQoJq8fW3iH = on0J0v1C0T4Vx5BAyNciCG <= xbDZHFjT9czSWoXqDrDalH; assign fWYsiC8varEjDaABQEOnHD = {L8G5zN2h3nNrCok5TCsJbE, rIIATJviRgNIQoJq8fW3iH}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : IcKFfaUrr3FW5eiYpHBh0G if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin jWzhv1CNrrkZ90yAhAoazF <= 14'b00000000000000; end else begin jWzhv1CNrrkZ90yAhAoazF <= fWYsiC8varEjDaABQEOnHD; end end assign m6rhgeyCXShlzRN5AMh18G = {DXqu7TpZsKBJkGAUCIfEdB, 2'b00}; assign GJygrD3xsfw2DPQ22BhMnF = (rIIATJviRgNIQoJq8fW3iH == 1'b0 ? m6rhgeyCXShlzRN5AMh18G : on0J0v1C0T4Vx5BAyNciCG); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : PebulLQF8uRrWOQ0S1MqbB if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin rqeR6AxGoUnIpcf8RFZE0C <= 28'b0000000000000000000000000000; end else begin rqeR6AxGoUnIpcf8RFZE0C <= GJygrD3xsfw2DPQ22BhMnF; end end assign uxJF4VESfR9zjMeGYtrIS = {rqeR6AxGoUnIpcf8RFZE0C, 2'b01}; assign a9YNARWK4HMkgu5zeMeFqB = {jWzhv1CNrrkZ90yAhAoazF, 2'b00}; assign OJCxI8u48szx5fkdxbfWjF = ({1'b0, uxJF4VESfR9zjMeGYtrIS}) + ({15'b0, a9YNARWK4HMkgu5zeMeFqB}); assign Nqy6crAgfKalgWwdaoPgWF = (OJCxI8u48szx5fkdxbfWjF[30] != 1'b0 ? 30'b111111111111111111111111111111 : OJCxI8u48szx5fkdxbfWjF[29:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : zijl3VQE0ZivHKrnknV0T if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin UVyVvhhWLxLhiHSNKkfKfE <= 32'b00000000000000000000000000000000; end else begin UVyVvhhWLxLhiHSNKkfKfE <= zjMYjjAxK45sdDEQ0XFXOG; end end assign VPMmTC28HmTVgoT6ZLk0CD = UVyVvhhWLxLhiHSNKkfKfE[31:2]; assign T4LoOhTfaEIFoiHehRN8gB = Nqy6crAgfKalgWwdaoPgWF <= VPMmTC28HmTVgoT6ZLk0CD; assign z7KS1tRTiUNV07mMLJEuKG = {jWzhv1CNrrkZ90yAhAoazF, T4LoOhTfaEIFoiHehRN8gB}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : r4sMtNTnn0C61Z9TeBBCEE if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin TKE1ENeioNod9UMhIzVfSH <= 15'b000000000000000; end else begin TKE1ENeioNod9UMhIzVfSH <= z7KS1tRTiUNV07mMLJEuKG; end end assign nkdnEk7YtJ3W7AmLNPDo = {rqeR6AxGoUnIpcf8RFZE0C, 2'b00}; assign y5KCvh2zjCyG1LFiVsUMYcD = (T4LoOhTfaEIFoiHehRN8gB == 1'b0 ? nkdnEk7YtJ3W7AmLNPDo : Nqy6crAgfKalgWwdaoPgWF); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : f9SedVstZyvPr0vo4Nl0pZF if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin cZ0D6qUE7QWbwvVcyFlvNC <= 30'b000000000000000000000000000000; end else begin cZ0D6qUE7QWbwvVcyFlvNC <= y5KCvh2zjCyG1LFiVsUMYcD; end end assign zD10HQPaWNtGjDTMJz3GSH = {cZ0D6qUE7QWbwvVcyFlvNC, 2'b01}; assign d9bLW3agjcpEpWrolrVdsmC = {TKE1ENeioNod9UMhIzVfSH, 2'b00}; assign QJOFvqfWKUFnEFOqoOrxWG = ({1'b0, zD10HQPaWNtGjDTMJz3GSH}) + ({16'b0, d9bLW3agjcpEpWrolrVdsmC}); assign z1qYldk164H9FNaPWpn6hF = (QJOFvqfWKUFnEFOqoOrxWG[32] != 1'b0 ? 32'b11111111111111111111111111111111 : QJOFvqfWKUFnEFOqoOrxWG[31:0]); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : PiQ9IEK7vsPtjrDsIFlXn if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin m47DvfSzOdN9OKy9YulLguB <= 32'b00000000000000000000000000000000; end else begin m47DvfSzOdN9OKy9YulLguB <= UVyVvhhWLxLhiHSNKkfKfE; end end assign cpmy5PzhVLGXdDoyCkUWiD = z1qYldk164H9FNaPWpn6hF <= m47DvfSzOdN9OKy9YulLguB; assign LPQDAvbrOjkrOtmk9vzPJB = {TKE1ENeioNod9UMhIzVfSH, cpmy5PzhVLGXdDoyCkUWiD}; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : ZhC3on7NcVQXKKMO6rEb9F if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin agalUIcyHoMvnBXt7uR1FE <= 16'b0000000000000000; end else begin agalUIcyHoMvnBXt7uR1FE <= LPQDAvbrOjkrOtmk9vzPJB; end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : l7YDg91XXtUA5EBaC0urXD if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin VDuk3ojf4kqPZHi2nVzzSD[0] <= 16'b0000000000000000; VDuk3ojf4kqPZHi2nVzzSD[1] <= 16'b0000000000000000; end else begin VDuk3ojf4kqPZHi2nVzzSD[0] <= xzmEHvAakc16M7C3TuYQlF[0]; VDuk3ojf4kqPZHi2nVzzSD[1] <= xzmEHvAakc16M7C3TuYQlF[1]; end end assign n6vRpiFqkFIHzpDYbJGYiD = VDuk3ojf4kqPZHi2nVzzSD[1]; assign xzmEHvAakc16M7C3TuYQlF[0] = agalUIcyHoMvnBXt7uR1FE; assign xzmEHvAakc16M7C3TuYQlF[1] = VDuk3ojf4kqPZHi2nVzzSD[0]; assign q3w3Ce5AlDM2h7wxTsVajWB = n6vRpiFqkFIHzpDYbJGYiD; assign s7ASYYS329kRVgP7KY37Y = q3w3Ce5AlDM2h7wxTsVajWB; endmodule