`timescale 1 ns / 1 ns module d4QD8esP7XdYbm4O3mpV7GH (v04pHKxyc2sPW047bbyUgE, JAMOfrNHxGSYDF0urqkLN, w3gGIVls9UktX3B50XtCM9D, PkjFB7tzez7RAWc2cSLnBD, cuDt5zGIRdJYB1ZsmaWyNE, a1hhzPnRvmngQQ69MdICU7C, PF6wwTYP1q9nJ5YwMDlzXE, NunEp0PDJBOuCyVdY3ejIC, zTC5dHloAQWrunmpBf9AuG, d8pq1PMmLZANfmOanWWlBYF, xj2txhdk3kH1ioK0rKOVrG, R6zf5iqRNVEGVBO8egq8kF, mdal5obekPJm0ao7ZiZ4cF, q4mhS1P9mOTwehAXXNmhxF, vyWRmDyKy2RVVIdRBtzV5F, SRoFC9yIIwEIUwYpoyy0QF, wpHiLzmis5ns3l38MddOzE, j963sPBld8mpm71sqcvb8WF, Ic4vfYy6jnxaw8uXI98INH, x2KkW4HKTQgVBmVskDu4RD, g1D8wSsV4Ksuy5G0qxKYMs); input v04pHKxyc2sPW047bbyUgE; input JAMOfrNHxGSYDF0urqkLN; input signed [15:0] w3gGIVls9UktX3B50XtCM9D; input signed [15:0] PkjFB7tzez7RAWc2cSLnBD; input signed [15:0] cuDt5zGIRdJYB1ZsmaWyNE; input signed [15:0] a1hhzPnRvmngQQ69MdICU7C; input signed [15:0] PF6wwTYP1q9nJ5YwMDlzXE; input signed [15:0] NunEp0PDJBOuCyVdY3ejIC; input signed [15:0] zTC5dHloAQWrunmpBf9AuG; input signed [15:0] d8pq1PMmLZANfmOanWWlBYF; input xj2txhdk3kH1ioK0rKOVrG; input R6zf5iqRNVEGVBO8egq8kF; output signed [15:0] mdal5obekPJm0ao7ZiZ4cF; output signed [15:0] q4mhS1P9mOTwehAXXNmhxF; output signed [15:0] vyWRmDyKy2RVVIdRBtzV5F; output signed [15:0] SRoFC9yIIwEIUwYpoyy0QF; output signed [15:0] wpHiLzmis5ns3l38MddOzE; output signed [15:0] j963sPBld8mpm71sqcvb8WF; output signed [15:0] Ic4vfYy6jnxaw8uXI98INH; output signed [15:0] x2KkW4HKTQgVBmVskDu4RD; output g1D8wSsV4Ksuy5G0qxKYMs; wire Ebx0yJLDGKevxkqzRPIfvG; wire signed [15:0] VZb9IGNA6knXVYHTLgj0yE; wire signed [15:0] GfOU8VnvrygAR1sS2nk8nB; wire signed [15:0] mf8WSHlMlZlNiovf5yywn; wire signed [15:0] qe6tQ6Jsl5fvHsen124cfC; wire Z7ZDy0EvwvoCh1zahAqvSF; wire signed [15:0] B58twvtfgVWGK5P29KavtH; wire signed [15:0] qhk6Uhwhppvpssqm7Nh6XE; wire signed [15:0] k3VfrgkD6DWITJL9WW5W4D; wire signed [15:0] pPn6MVGqBLqJ0xzN2WYfFG; wire jNZ4xylBKAANfCL11XNxzB; wire signed [15:0] BpNlQ4LQUlVTEBlULLLjXE; wire signed [15:0] TlwXorPjcpNngmZL5m6lQG; wire signed [15:0] v67zkeDCrQzNzBtQlbUWdG; wire signed [15:0] OIn98Mhn9PlHJx0jNKukHB; wire signed [15:0] VWSiqDgxQN9a2J7zRy3p4E; wire signed [15:0] LhqlKpPzANkuN2xC8HYciC; wire signed [15:0] OUMqBzkN19EDa2VTABMa2E; wire signed [15:0] qbEnMIxMUsx8pYkF1gFd7D; wire signed [15:0] A5SQIaNgqW7DcTqQkKRVeD; wire signed [15:0] GaetbCaMty7UkzjqNoYErC; wire signed [15:0] M5AqS9R7rFTkWxwo8io2rH; wire signed [15:0] lcJo4MnEaj41ofRAtLkn4D; wire Pq4nKEqqr18aLXK1kX1dfH; reg signed [15:0] XQltXNYzwWy18SM8pDhf8 [0:2]; wire signed [15:0] V1YnWmj1nZzru97DWQqYdE [0:2]; wire signed [15:0] FPJLoZTbR5NUHIeb5WjctB; reg signed [15:0] TqWcgwsoO3Igmoq6nH36SB [0:2]; wire signed [15:0] pIqvCE2ZCwGFIfCd4j88bF [0:2]; wire signed [15:0] j7QbZWviLec2smu8yuKCIPF; reg [0:2] c5tyBuJoNrswqnLWL1VV0SB; wire [0:2] mqwYm78twnDBgE5C13tVbH; wire pCWATI9lTIGbmXTtLuLAGB; wire signed [15:0] zFuIFDmench8v1O4yXu4jG; wire signed [15:0] dQK1re9uLGxG0WuVGLoXdH; wire kIsHJAwQMWbIiCsXfX1rTG; wire yTf5WZbZOLm2uKwJmXk5sG; wire wGlnEfCkRPxniOjCaZH6XG; wire RDvlVEJspE7WkJvNmR8a6C; wire signed [15:0] H8Iagd3fwKKnwcTjUyOkqB; wire signed [15:0] CVOHwOszKLN4rogfAKlMXB; wire DZol1WsbVnSldsei0SiI9E; wire sIaC8spfzCmUwexq8stmB; wire zqdZMmoxIs9zmnL4kATVuC; wire a8rK4qdEuNCWHLdYbR2f8; wire O6TgnxqnGk692qEmnZQFTC; wire XfCDnggI1Y1qaMzSOLL0TD; wire signed [15:0] qfBqSs1n7vrUenPHRhvA4E; wire signed [15:0] s1Ni5BKBwo5acvXPnlIkC4D; wire NMWfejbHi1tIjFkylFWDkC; reg signed [15:0] LqbGk6Fit5FCOuam4sOAAD [0:2]; wire signed [15:0] Bi3HF1UTdSkQGHjQ4xRwvF [0:2]; wire signed [15:0] lyOqtmFbWBeDZLo4tO89VD; reg signed [15:0] yLZlCsGdKifpjAYDy4DDED [0:2]; wire signed [15:0] o2lMuceP2Zz2x444DyOgERH [0:2]; wire signed [15:0] nMEIHp8iZdLbxWoHks1NAB; reg [0:2] KyQ2PfyWtleyBDhGs5a1gF; wire [0:2] l750CVLudfD6Rvkr3byjjvH; wire v6PtMRDEb2KzMpzXWCSiwkB; wire signed [15:0] HXT3YNFExOHI94Xq9VVUBG; wire signed [15:0] EI1r2DTkmcgS5siR9DUFpG; wire NHkD6RGVcC6B7ibmcHypOC; wire [1:0] u6oVvmCf0f079jLPodlV5B; wire qv4pS1KBm1VYTuOTZHo04F; wire LSv5mOYTPLq5vaIpiVTypC; wire signed [15:0] zsayMT6gR21wpeAixbNYEF; wire signed [15:0] CaTCMDu7mVwW7eYB1tjZ5; wire Ck459KQ1C8vRbine3lrkt; wire DCqZJgzh8RI4wgf1TYRoc; wire [2:0] MCqIdNMOB0Mg1cefHLMjpH; wire j41GwwL8b9NI9l6ZScQ1PbG; wire i8H7HzN3cvjFks6MZ5qaqF; wire SAcShGLK2YZQrWHGqGVvjD; wire signed [15:0] rFr1ZhZNiURIbPFlZaI4kB; wire signed [15:0] gJidztDROiWi1BoJ2KzqKB; wire mm30CTneMiOZJcmmoHkb2D; reg signed [15:0] cVMiV2j8qD0P3CVc315hn [0:2]; wire signed [15:0] a9iZ9svlbzlFdVAGUFPTY [0:2]; wire signed [15:0] HeHFnbPrPBgeQHatNQHc0; reg signed [15:0] u2yic2bBqAL2jFtl9bgNqD [0:2]; wire signed [15:0] rKHf7GW9kd2HwW2mmfwvqC [0:2]; wire signed [15:0] gGCeJXlbwaFahBmsH6mMkF; reg [0:2] qM3kFDhftMVWrl1HT1qB4F; wire [0:2] eHbdLpdf2r0lFYM9BhuRoB; wire l9QVSAqS6jsMaipvGnosLD; wire signed [15:0] xj58yogg0Lfx8mMLdFuZsE; wire signed [15:0] IGbVPdIVOky0HoXMmdGGQH; wire wf5f4XnltnQYt1bEDWEp0F; reg VzGh5mviLsfsu1Hv3n1l5C; wire FUS5RSCs5VyI8J3rzh0AIE; wire [3:0] g1oJwDFAtNAcPvLahTlMEB; wire Q7D2KKVRLkwEPktPhyCkSD; wire signed [15:0] g1qVkXUxL7Fv5Vq7GJfmGVG; wire signed [15:0] UAWBm55LOUyC0bgEaA5EMC; wire g3JMyJIWtKhpmOxBRsFzIOH; wire j8MMagsoA5t6IysA2ZD3X4F; wire signed [15:0] aydyoHsGbz0wVGlm34qlsB; wire signed [15:0] H0BpAwmwCivCDsbLQ5qvCC; wire signed [15:0] s1N0USypDrc4xyzxc4XEMr; wire signed [15:0] sZ7bCwrhIAA80IOhzh695; reg signed [15:0] f69xGE65xXz2LbsT91hgR8G [0:2]; wire signed [15:0] v4gfbuVl5KUcQzK24qqOvB [0:2]; wire signed [15:0] DbYwoM2JCYD9mwcRRKmb6G; reg signed [15:0] v2G3ZeHqmqPQjfLNmkS0OrG [0:2]; wire signed [15:0] BrQqlwQZdOtmNiJOrBili [0:2]; wire signed [15:0] WbySmFpEqdJe6nrpd6KgG; wire signed [15:0] i4y6Td18s9Zr0JbepLQtjC; wire signed [15:0] k3FlrGNoOUOhUgHDIDYGouE; wire signed [15:0] t30W3eeadZl9O9RnQCafyED; wire signed [15:0] flGpcmOyc38fKmqiV5eQvF; wire signed [15:0] CBqrXFTnHQDD2JNQjTxpkH; wire signed [15:0] dYQ3fSOENqw4ZimOQmMMTH; reg signed [15:0] k11T3BX1fbEFyiI1W12X7 [0:2]; wire signed [15:0] VpKk1YVVYHSJ6RsO9pshiB [0:2]; wire signed [15:0] lSTAIQPANZYVi9u1bQJbfC; reg signed [15:0] RAKTymlGVAtDEhqm1mBWKC [0:2]; wire signed [15:0] yyMRtRepkZFuqH6zjb0hbC [0:2]; wire signed [15:0] hh7M8p6TyfjHKgE0YxcN3; wire signed [15:0] FB6nKajjqrTT1538hBpQ9C; wire signed [15:0] XcmpMS0nhYnUzTPGBkEmmF; wire signed [15:0] OAkG388GVoqfAFfrsC3Z3; wire signed [15:0] DP58bSOk4VSBFH6tnqlVTH; wire signed [15:0] oEtRmwXRZkMV2JHZdumYM; wire signed [15:0] ABAJKgUy1j1LH4rwhRtEnG; reg signed [15:0] k9BY0fd7LFxuaZBtnq2NstC [0:2]; wire signed [15:0] mTZgUkGw3710r8TqEV6XWF [0:2]; wire signed [15:0] PLuy3wDbVIiPXXOVcF7GXC; reg signed [15:0] k8gGlV5iKkuIBPqjsMS5KF [0:2]; wire signed [15:0] jVudy6rBy3pL4AAajihjvH [0:2]; wire signed [15:0] wt5uyiFelHvOxXII8I6cTH; wire signed [15:0] gQ8ol00XUcRCyi5uaxpHDB; wire signed [15:0] rj0jYY5GSDAuDuCDoIpZ9C; wire signed [15:0] jZwXcJxnQcGGzLJPOScVqE; wire signed [15:0] hP5DBuEisrqC9fZ23jziMF; reg signed [15:0] x9EdsEkQtjpM4w517iGHzC [0:2]; wire signed [15:0] tnuZKwedoQlWAtzBo6aIZB [0:2]; wire signed [15:0] risZnLFYvPBrH1cy6dfHMF; reg signed [15:0] KmuHj4FutgT59Q7oCiggpD [0:2]; wire signed [15:0] UFFCUGMTW5jYs8JEV3j3KC [0:2]; wire signed [15:0] y3mUIhc5hpdbI6gB0Klf3MH; wire signed [15:0] UlGc2PVtJa9BNobxUHDxSG; wire signed [15:0] pdTCH0gTlgy9qR74rtvuBE; wire signed [15:0] msLJn85q5aDnigXPSLnA9F; wire signed [15:0] s8tbEDkTdSLkOXc5hVDArH; wire signed [15:0] ACHpp43jQbQJO4HdGlLQ0B; wire signed [15:0] BJNXQzaMpa7r8LYTHlOrBD; reg signed [15:0] appAG8sqUT59wY8ObKEssF [0:2]; wire signed [15:0] d21AAbScpxqwLWzuGxj8ajB [0:2]; wire signed [15:0] BXAaMHpKzPpYZGFRqoevNE; reg signed [15:0] pISZVQJtPY1M87J4LAx1MB [0:2]; wire signed [15:0] EwyTeOtw0Znxv6WUZIsKtH [0:2]; wire signed [15:0] czP63K90EaJdtsY9EHZ30D; wire signed [15:0] mxtJaiWQH83FcZ66WqnMiH; wire signed [15:0] MtlWbaE0z2xTCIy368PlWF; wire signed [15:0] Sek0doTmbyRuabtHW5JKgH; wire signed [15:0] h4q2yYljVPy2UhMxEpHXfqG; wire signed [15:0] Ni5CWVNOepdNWeLhPbktyC; wire signed [15:0] oC9IZ8suhbNZiMMpUwYFZE; reg signed [15:0] ufyCKBsm7ZcDMoHa9lVT8B [0:2]; wire signed [15:0] lc0FzXjU6ruJOOuwpT5PQ [0:2]; wire signed [15:0] z6SwcDGEsoURdwbnSfOpHB; reg signed [15:0] f6n0j0rIhtlF1cK7ntOhdG [0:2]; wire signed [15:0] f8PGb7nqRvYgidEKAnbVYCF [0:2]; wire signed [15:0] pGKHaOZvJloUuxOXANTYZE; wire signed [15:0] feyfHDrrhsk9bdeB57O2c; wire signed [15:0] r2IKtvrSH76nVotfMIojNdD; wire signed [15:0] SmUoeWULdUSlbsjccscXpG; wire signed [15:0] qrJeNpaPfOy0pMCu40c1ME; reg signed [15:0] hDe4KgCGLUE2lc3mBRHUGE [0:2]; wire signed [15:0] ZvqDLDMtFPbHpUtzihpbXF [0:2]; wire signed [15:0] EiKTmNA9gqnqt6QU2ytsGF; reg signed [15:0] I3TwcvTY4hEZBUKyNKGQYH [0:2]; wire signed [15:0] ltutKZEJ3uAsYBtveZfxN [0:2]; wire signed [15:0] i0padod73DFvzROjA4fS2o; wire signed [15:0] mvb8xVo6CcFPFyQu3ctDE; wire signed [15:0] gC05dypmmuscVux3EfDHCD; wire signed [15:0] DxKKPTJNNNGcVbnDyBefdC; wire signed [15:0] z5IVnN9scVD1jMboeUZaZG; wire signed [15:0] y2F62Qir2uvIcDNjqoCgbPG; wire signed [15:0] eJSHu1mAvW9BzbMy0ufWWD; reg signed [15:0] h41dWYc0X3ZAsDk44FMtsTD [0:2]; wire signed [15:0] kZIaatjtNR5S1owTPfmSI [0:2]; wire signed [15:0] SNl44VPeKmo2uIh5zCljYE; reg signed [15:0] UbhppxZFtuRiGSMYxgMT2F [0:2]; wire signed [15:0] rk6XtqxIQmYnoKIvpO9PNH [0:2]; wire signed [15:0] AXkTVaeFKW3Cvod76gwXK; wire signed [15:0] PV2GPYF9MTfm6A3VIE3yL; wire signed [15:0] VMMfdu9AIUdQe4XcwZLbSC; wire signed [15:0] BSA6wYLjrd40iGAxWAWPUG; wire signed [15:0] mVsThSJWeEPGLaZQZJ476C; wire signed [15:0] Qjop49qrCNJ2RVI1tmxWK; wire signed [15:0] qtlf3VUxsnDXMsfKMVqqRD; reg signed [15:0] TGSVeodh4aSh5YMUFsJBpF [0:2]; wire signed [15:0] pKwMCjbBuwX4wlYrJtZeqH [0:2]; wire signed [15:0] T6wR1FRvpbz8HFANbQ6odH; reg signed [15:0] t1XxIWfdmuGYgMJ14AA5aoF [0:2]; wire signed [15:0] Ed8ZUSDNSkOaxlQSyerJMG [0:2]; wire signed [15:0] c88iPPDCYH3uMXl21XZoi8D; wire signed [15:0] RRE1h6KsUsyxLABwNoPOPB; wire signed [15:0] vM9w9urjKvIy07zqFkMIPF; wire signed [15:0] tZCSNlfV8pGx0wl9RXazqC; wire signed [15:0] vuJEKfnV5iqg56DSJMMzfH; wire ICbriSzMXIBZ11lqkoCXnD; assign Ebx0yJLDGKevxkqzRPIfvG = 1'b0; assign VZb9IGNA6knXVYHTLgj0yE = w3gGIVls9UktX3B50XtCM9D; assign GfOU8VnvrygAR1sS2nk8nB = PF6wwTYP1q9nJ5YwMDlzXE; assign mf8WSHlMlZlNiovf5yywn = PkjFB7tzez7RAWc2cSLnBD; assign qe6tQ6Jsl5fvHsen124cfC = NunEp0PDJBOuCyVdY3ejIC; assign Z7ZDy0EvwvoCh1zahAqvSF = (xj2txhdk3kH1ioK0rKOVrG != 1'b0 ? 1'b1 : 1'b0); n18IkTlDKVWTnppeBlI84nG u4hlhjEy5S0jdWbgdAzINDD (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .EnlAo7K66kKuzHIKWLmc1F(VZb9IGNA6knXVYHTLgj0yE), .ew3EeLap6s8rXmNrsqaTWH(GfOU8VnvrygAR1sS2nk8nB), .IPh1M0O3x0ioGlon72MROG(mf8WSHlMlZlNiovf5yywn), .Mt05SNCQbo0cCPNa1yEFyF(qe6tQ6Jsl5fvHsen124cfC), .Z7ZDy0EvwvoCh1zahAqvSF(Z7ZDy0EvwvoCh1zahAqvSF), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .B58twvtfgVWGK5P29KavtH(B58twvtfgVWGK5P29KavtH), .qhk6Uhwhppvpssqm7Nh6XE(qhk6Uhwhppvpssqm7Nh6XE), .k3VfrgkD6DWITJL9WW5W4D(k3VfrgkD6DWITJL9WW5W4D), .pPn6MVGqBLqJ0xzN2WYfFG(pPn6MVGqBLqJ0xzN2WYfFG), .jNZ4xylBKAANfCL11XNxzB(jNZ4xylBKAANfCL11XNxzB) ); assign BpNlQ4LQUlVTEBlULLLjXE = cuDt5zGIRdJYB1ZsmaWyNE; assign TlwXorPjcpNngmZL5m6lQG = zTC5dHloAQWrunmpBf9AuG; assign v67zkeDCrQzNzBtQlbUWdG = a1hhzPnRvmngQQ69MdICU7C; assign OIn98Mhn9PlHJx0jNKukHB = d8pq1PMmLZANfmOanWWlBYF; GpUftF8ITUnSwAZhyOk5qD KLMaXcYHHyApMQQHB9ZGnC (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .qmhLAZZAHFrO09l1zXnPRC(BpNlQ4LQUlVTEBlULLLjXE), .JMtgCMT5TVzyJSn9uILA1(TlwXorPjcpNngmZL5m6lQG), .xYJCS7zMCKI1yYR3Bx1XrD(v67zkeDCrQzNzBtQlbUWdG), .AaqUpSvCGAV1YR86nIsLWH(OIn98Mhn9PlHJx0jNKukHB), .Z7ZDy0EvwvoCh1zahAqvSF(Z7ZDy0EvwvoCh1zahAqvSF), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .VWSiqDgxQN9a2J7zRy3p4E(VWSiqDgxQN9a2J7zRy3p4E), .LhqlKpPzANkuN2xC8HYciC(LhqlKpPzANkuN2xC8HYciC), .OUMqBzkN19EDa2VTABMa2E(OUMqBzkN19EDa2VTABMa2E), .qbEnMIxMUsx8pYkF1gFd7D(qbEnMIxMUsx8pYkF1gFd7D) ); xRgm1KQSpBEMURvTRAnYsB lm0pV74Hf3yaqeAtQU1kHF (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .Ebx0yJLDGKevxkqzRPIfvG(Ebx0yJLDGKevxkqzRPIfvG), .B58twvtfgVWGK5P29KavtH(B58twvtfgVWGK5P29KavtH), .qhk6Uhwhppvpssqm7Nh6XE(qhk6Uhwhppvpssqm7Nh6XE), .VWSiqDgxQN9a2J7zRy3p4E(VWSiqDgxQN9a2J7zRy3p4E), .LhqlKpPzANkuN2xC8HYciC(LhqlKpPzANkuN2xC8HYciC), .jNZ4xylBKAANfCL11XNxzB(jNZ4xylBKAANfCL11XNxzB), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .A5SQIaNgqW7DcTqQkKRVeD(A5SQIaNgqW7DcTqQkKRVeD), .GaetbCaMty7UkzjqNoYErC(GaetbCaMty7UkzjqNoYErC), .k3VfrgkD6DWITJL9WW5W4D(M5AqS9R7rFTkWxwo8io2rH), .pPn6MVGqBLqJ0xzN2WYfFG(lcJo4MnEaj41ofRAtLkn4D), .Pq4nKEqqr18aLXK1kX1dfH(Pq4nKEqqr18aLXK1kX1dfH) ); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : MczQYJ6MT1pYZD7C1UhQv if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin XQltXNYzwWy18SM8pDhf8[0] <= 16'sb0000000000000000; XQltXNYzwWy18SM8pDhf8[1] <= 16'sb0000000000000000; XQltXNYzwWy18SM8pDhf8[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin XQltXNYzwWy18SM8pDhf8[0] <= 16'sb0000000000000000; XQltXNYzwWy18SM8pDhf8[1] <= 16'sb0000000000000000; XQltXNYzwWy18SM8pDhf8[2] <= 16'sb0000000000000000; end else begin XQltXNYzwWy18SM8pDhf8[0] <= V1YnWmj1nZzru97DWQqYdE[0]; XQltXNYzwWy18SM8pDhf8[1] <= V1YnWmj1nZzru97DWQqYdE[1]; XQltXNYzwWy18SM8pDhf8[2] <= V1YnWmj1nZzru97DWQqYdE[2]; end end end assign FPJLoZTbR5NUHIeb5WjctB = XQltXNYzwWy18SM8pDhf8[2]; assign V1YnWmj1nZzru97DWQqYdE[0] = A5SQIaNgqW7DcTqQkKRVeD; assign V1YnWmj1nZzru97DWQqYdE[1] = XQltXNYzwWy18SM8pDhf8[0]; assign V1YnWmj1nZzru97DWQqYdE[2] = XQltXNYzwWy18SM8pDhf8[1]; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : xwyxj2YIc64Lxvl4r8S8mG if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin TqWcgwsoO3Igmoq6nH36SB[0] <= 16'sb0000000000000000; TqWcgwsoO3Igmoq6nH36SB[1] <= 16'sb0000000000000000; TqWcgwsoO3Igmoq6nH36SB[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin TqWcgwsoO3Igmoq6nH36SB[0] <= 16'sb0000000000000000; TqWcgwsoO3Igmoq6nH36SB[1] <= 16'sb0000000000000000; TqWcgwsoO3Igmoq6nH36SB[2] <= 16'sb0000000000000000; end else begin TqWcgwsoO3Igmoq6nH36SB[0] <= pIqvCE2ZCwGFIfCd4j88bF[0]; TqWcgwsoO3Igmoq6nH36SB[1] <= pIqvCE2ZCwGFIfCd4j88bF[1]; TqWcgwsoO3Igmoq6nH36SB[2] <= pIqvCE2ZCwGFIfCd4j88bF[2]; end end end assign j7QbZWviLec2smu8yuKCIPF = TqWcgwsoO3Igmoq6nH36SB[2]; assign pIqvCE2ZCwGFIfCd4j88bF[0] = GaetbCaMty7UkzjqNoYErC; assign pIqvCE2ZCwGFIfCd4j88bF[1] = TqWcgwsoO3Igmoq6nH36SB[0]; assign pIqvCE2ZCwGFIfCd4j88bF[2] = TqWcgwsoO3Igmoq6nH36SB[1]; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : L1HBH8O5DRbGBa9XvBX70C if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin c5tyBuJoNrswqnLWL1VV0SB[0] <= 1'b0; c5tyBuJoNrswqnLWL1VV0SB[1] <= 1'b0; c5tyBuJoNrswqnLWL1VV0SB[2] <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin c5tyBuJoNrswqnLWL1VV0SB[0] <= 1'b0; c5tyBuJoNrswqnLWL1VV0SB[1] <= 1'b0; c5tyBuJoNrswqnLWL1VV0SB[2] <= 1'b0; end else begin c5tyBuJoNrswqnLWL1VV0SB[0] <= mqwYm78twnDBgE5C13tVbH[0]; c5tyBuJoNrswqnLWL1VV0SB[1] <= mqwYm78twnDBgE5C13tVbH[1]; c5tyBuJoNrswqnLWL1VV0SB[2] <= mqwYm78twnDBgE5C13tVbH[2]; end end end assign pCWATI9lTIGbmXTtLuLAGB = c5tyBuJoNrswqnLWL1VV0SB[2]; assign mqwYm78twnDBgE5C13tVbH[0] = Pq4nKEqqr18aLXK1kX1dfH; assign mqwYm78twnDBgE5C13tVbH[1] = c5tyBuJoNrswqnLWL1VV0SB[0]; assign mqwYm78twnDBgE5C13tVbH[2] = c5tyBuJoNrswqnLWL1VV0SB[1]; t3fQLgkwcS9J9XUJPuAx7jC qTfyhdbQzAKcKbDpRJj8yG (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .Pq4nKEqqr18aLXK1kX1dfH(Pq4nKEqqr18aLXK1kX1dfH), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .zFuIFDmench8v1O4yXu4jG(zFuIFDmench8v1O4yXu4jG), .dQK1re9uLGxG0WuVGLoXdH(dQK1re9uLGxG0WuVGLoXdH) ); c5frKpr1OF9l0qPiwsMhI2 JSNmXQ0YI7nAzGfsGLG1UC (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .kIsHJAwQMWbIiCsXfX1rTG(kIsHJAwQMWbIiCsXfX1rTG), .DKGIysOp4cb2Wy4ifYHB8D(kIsHJAwQMWbIiCsXfX1rTG), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .yTf5WZbZOLm2uKwJmXk5sG(yTf5WZbZOLm2uKwJmXk5sG), .wGlnEfCkRPxniOjCaZH6XG(wGlnEfCkRPxniOjCaZH6XG), .RDvlVEJspE7WkJvNmR8a6C(RDvlVEJspE7WkJvNmR8a6C) ); OwsLDamo9WkovW7t04kXBG rKXyl8hgTMym1rEDLsJaOB (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .FPJLoZTbR5NUHIeb5WjctB(FPJLoZTbR5NUHIeb5WjctB), .j7QbZWviLec2smu8yuKCIPF(j7QbZWviLec2smu8yuKCIPF), .pCWATI9lTIGbmXTtLuLAGB(pCWATI9lTIGbmXTtLuLAGB), .yTf5WZbZOLm2uKwJmXk5sG(yTf5WZbZOLm2uKwJmXk5sG), .wGlnEfCkRPxniOjCaZH6XG(wGlnEfCkRPxniOjCaZH6XG), .zFuIFDmench8v1O4yXu4jG(zFuIFDmench8v1O4yXu4jG), .dQK1re9uLGxG0WuVGLoXdH(dQK1re9uLGxG0WuVGLoXdH), .RDvlVEJspE7WkJvNmR8a6C(RDvlVEJspE7WkJvNmR8a6C), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .H8Iagd3fwKKnwcTjUyOkqB(H8Iagd3fwKKnwcTjUyOkqB), .CVOHwOszKLN4rogfAKlMXB(CVOHwOszKLN4rogfAKlMXB), .DZol1WsbVnSldsei0SiI9E(DZol1WsbVnSldsei0SiI9E), .kIsHJAwQMWbIiCsXfX1rTG(kIsHJAwQMWbIiCsXfX1rTG) ); m0wR0p8t3oV06dM5Osycg9 z962IOrouyDUWLniu10oD3C (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .DZol1WsbVnSldsei0SiI9E(DZol1WsbVnSldsei0SiI9E), .sIaC8spfzCmUwexq8stmB(sIaC8spfzCmUwexq8stmB), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .zqdZMmoxIs9zmnL4kATVuC(zqdZMmoxIs9zmnL4kATVuC), .a8rK4qdEuNCWHLdYbR2f8(a8rK4qdEuNCWHLdYbR2f8), .O6TgnxqnGk692qEmnZQFTC(O6TgnxqnGk692qEmnZQFTC), .XfCDnggI1Y1qaMzSOLL0TD(XfCDnggI1Y1qaMzSOLL0TD) ); iUXDhKLNoaXRbJ8f5ydmRD onkga9gnAWHYkWnfgU4ydB (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .H8Iagd3fwKKnwcTjUyOkqB(H8Iagd3fwKKnwcTjUyOkqB), .CVOHwOszKLN4rogfAKlMXB(CVOHwOszKLN4rogfAKlMXB), .DZol1WsbVnSldsei0SiI9E(DZol1WsbVnSldsei0SiI9E), .zqdZMmoxIs9zmnL4kATVuC(zqdZMmoxIs9zmnL4kATVuC), .a8rK4qdEuNCWHLdYbR2f8(a8rK4qdEuNCWHLdYbR2f8), .O6TgnxqnGk692qEmnZQFTC(O6TgnxqnGk692qEmnZQFTC), .XfCDnggI1Y1qaMzSOLL0TD(XfCDnggI1Y1qaMzSOLL0TD), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .qfBqSs1n7vrUenPHRhvA4E(qfBqSs1n7vrUenPHRhvA4E), .s1Ni5BKBwo5acvXPnlIkC4D(s1Ni5BKBwo5acvXPnlIkC4D), .NMWfejbHi1tIjFkylFWDkC(NMWfejbHi1tIjFkylFWDkC), .sIaC8spfzCmUwexq8stmB(sIaC8spfzCmUwexq8stmB) ); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : s2CWr6rrksK4W7N0omU97HD if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin LqbGk6Fit5FCOuam4sOAAD[0] <= 16'sb0000000000000000; LqbGk6Fit5FCOuam4sOAAD[1] <= 16'sb0000000000000000; LqbGk6Fit5FCOuam4sOAAD[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin LqbGk6Fit5FCOuam4sOAAD[0] <= 16'sb0000000000000000; LqbGk6Fit5FCOuam4sOAAD[1] <= 16'sb0000000000000000; LqbGk6Fit5FCOuam4sOAAD[2] <= 16'sb0000000000000000; end else begin LqbGk6Fit5FCOuam4sOAAD[0] <= Bi3HF1UTdSkQGHjQ4xRwvF[0]; LqbGk6Fit5FCOuam4sOAAD[1] <= Bi3HF1UTdSkQGHjQ4xRwvF[1]; LqbGk6Fit5FCOuam4sOAAD[2] <= Bi3HF1UTdSkQGHjQ4xRwvF[2]; end end end assign lyOqtmFbWBeDZLo4tO89VD = LqbGk6Fit5FCOuam4sOAAD[2]; assign Bi3HF1UTdSkQGHjQ4xRwvF[0] = qfBqSs1n7vrUenPHRhvA4E; assign Bi3HF1UTdSkQGHjQ4xRwvF[1] = LqbGk6Fit5FCOuam4sOAAD[0]; assign Bi3HF1UTdSkQGHjQ4xRwvF[2] = LqbGk6Fit5FCOuam4sOAAD[1]; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : k1Zsi6BUVrSUjLbIYwh26G if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin yLZlCsGdKifpjAYDy4DDED[0] <= 16'sb0000000000000000; yLZlCsGdKifpjAYDy4DDED[1] <= 16'sb0000000000000000; yLZlCsGdKifpjAYDy4DDED[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin yLZlCsGdKifpjAYDy4DDED[0] <= 16'sb0000000000000000; yLZlCsGdKifpjAYDy4DDED[1] <= 16'sb0000000000000000; yLZlCsGdKifpjAYDy4DDED[2] <= 16'sb0000000000000000; end else begin yLZlCsGdKifpjAYDy4DDED[0] <= o2lMuceP2Zz2x444DyOgERH[0]; yLZlCsGdKifpjAYDy4DDED[1] <= o2lMuceP2Zz2x444DyOgERH[1]; yLZlCsGdKifpjAYDy4DDED[2] <= o2lMuceP2Zz2x444DyOgERH[2]; end end end assign nMEIHp8iZdLbxWoHks1NAB = yLZlCsGdKifpjAYDy4DDED[2]; assign o2lMuceP2Zz2x444DyOgERH[0] = s1Ni5BKBwo5acvXPnlIkC4D; assign o2lMuceP2Zz2x444DyOgERH[1] = yLZlCsGdKifpjAYDy4DDED[0]; assign o2lMuceP2Zz2x444DyOgERH[2] = yLZlCsGdKifpjAYDy4DDED[1]; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : TPi3Fu9uFLztbkFwa0H53D if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin KyQ2PfyWtleyBDhGs5a1gF[0] <= 1'b0; KyQ2PfyWtleyBDhGs5a1gF[1] <= 1'b0; KyQ2PfyWtleyBDhGs5a1gF[2] <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin KyQ2PfyWtleyBDhGs5a1gF[0] <= 1'b0; KyQ2PfyWtleyBDhGs5a1gF[1] <= 1'b0; KyQ2PfyWtleyBDhGs5a1gF[2] <= 1'b0; end else begin KyQ2PfyWtleyBDhGs5a1gF[0] <= l750CVLudfD6Rvkr3byjjvH[0]; KyQ2PfyWtleyBDhGs5a1gF[1] <= l750CVLudfD6Rvkr3byjjvH[1]; KyQ2PfyWtleyBDhGs5a1gF[2] <= l750CVLudfD6Rvkr3byjjvH[2]; end end end assign v6PtMRDEb2KzMpzXWCSiwkB = KyQ2PfyWtleyBDhGs5a1gF[2]; assign l750CVLudfD6Rvkr3byjjvH[0] = NMWfejbHi1tIjFkylFWDkC; assign l750CVLudfD6Rvkr3byjjvH[1] = KyQ2PfyWtleyBDhGs5a1gF[0]; assign l750CVLudfD6Rvkr3byjjvH[2] = KyQ2PfyWtleyBDhGs5a1gF[1]; o3WOD3rXumRGZuWbQyHSTC mYbRzIp6fh5UU50NIPMlqE (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .NMWfejbHi1tIjFkylFWDkC(NMWfejbHi1tIjFkylFWDkC), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .HXT3YNFExOHI94Xq9VVUBG(HXT3YNFExOHI94Xq9VVUBG), .EI1r2DTkmcgS5siR9DUFpG(EI1r2DTkmcgS5siR9DUFpG) ); HMcgSDBQI8srN5Fet9wEnG K59tEegFJMrdmJIuWBI7q (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .NHkD6RGVcC6B7ibmcHypOC(NHkD6RGVcC6B7ibmcHypOC), .n6CG7K4rgMGw86VJoKnfuOD(NHkD6RGVcC6B7ibmcHypOC), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .u6oVvmCf0f079jLPodlV5B(u6oVvmCf0f079jLPodlV5B), .qv4pS1KBm1VYTuOTZHo04F(qv4pS1KBm1VYTuOTZHo04F), .LSv5mOYTPLq5vaIpiVTypC(LSv5mOYTPLq5vaIpiVTypC) ); y3RjWI2gAkcor9IfmoDAhWC YGfiJxj5wy9c9fxm8qBmQC (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .lyOqtmFbWBeDZLo4tO89VD(lyOqtmFbWBeDZLo4tO89VD), .nMEIHp8iZdLbxWoHks1NAB(nMEIHp8iZdLbxWoHks1NAB), .v6PtMRDEb2KzMpzXWCSiwkB(v6PtMRDEb2KzMpzXWCSiwkB), .u6oVvmCf0f079jLPodlV5B(u6oVvmCf0f079jLPodlV5B), .qv4pS1KBm1VYTuOTZHo04F(qv4pS1KBm1VYTuOTZHo04F), .HXT3YNFExOHI94Xq9VVUBG(HXT3YNFExOHI94Xq9VVUBG), .EI1r2DTkmcgS5siR9DUFpG(EI1r2DTkmcgS5siR9DUFpG), .LSv5mOYTPLq5vaIpiVTypC(LSv5mOYTPLq5vaIpiVTypC), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .zsayMT6gR21wpeAixbNYEF(zsayMT6gR21wpeAixbNYEF), .CaTCMDu7mVwW7eYB1tjZ5(CaTCMDu7mVwW7eYB1tjZ5), .Ck459KQ1C8vRbine3lrkt(Ck459KQ1C8vRbine3lrkt), .NHkD6RGVcC6B7ibmcHypOC(NHkD6RGVcC6B7ibmcHypOC) ); QNagGs9mRrlwXRNR72KVyF BoxmA9gUrcoGKTr1WWdljB (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .Ck459KQ1C8vRbine3lrkt(Ck459KQ1C8vRbine3lrkt), .DCqZJgzh8RI4wgf1TYRoc(DCqZJgzh8RI4wgf1TYRoc), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .MCqIdNMOB0Mg1cefHLMjpH(MCqIdNMOB0Mg1cefHLMjpH), .j41GwwL8b9NI9l6ZScQ1PbG(j41GwwL8b9NI9l6ZScQ1PbG), .i8H7HzN3cvjFks6MZ5qaqF(i8H7HzN3cvjFks6MZ5qaqF), .SAcShGLK2YZQrWHGqGVvjD(SAcShGLK2YZQrWHGqGVvjD) ); AvW45ZD2J4hIv4kcbbeCqF v4tQ5NbkvrLEoEVGS2hwT8F (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .zsayMT6gR21wpeAixbNYEF(zsayMT6gR21wpeAixbNYEF), .CaTCMDu7mVwW7eYB1tjZ5(CaTCMDu7mVwW7eYB1tjZ5), .Ck459KQ1C8vRbine3lrkt(Ck459KQ1C8vRbine3lrkt), .MCqIdNMOB0Mg1cefHLMjpH(MCqIdNMOB0Mg1cefHLMjpH), .j41GwwL8b9NI9l6ZScQ1PbG(j41GwwL8b9NI9l6ZScQ1PbG), .i8H7HzN3cvjFks6MZ5qaqF(i8H7HzN3cvjFks6MZ5qaqF), .SAcShGLK2YZQrWHGqGVvjD(SAcShGLK2YZQrWHGqGVvjD), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .rFr1ZhZNiURIbPFlZaI4kB(rFr1ZhZNiURIbPFlZaI4kB), .gJidztDROiWi1BoJ2KzqKB(gJidztDROiWi1BoJ2KzqKB), .mm30CTneMiOZJcmmoHkb2D(mm30CTneMiOZJcmmoHkb2D), .DCqZJgzh8RI4wgf1TYRoc(DCqZJgzh8RI4wgf1TYRoc) ); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : IBmSJmjQmOQZECy1AykU1D if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin cVMiV2j8qD0P3CVc315hn[0] <= 16'sb0000000000000000; cVMiV2j8qD0P3CVc315hn[1] <= 16'sb0000000000000000; cVMiV2j8qD0P3CVc315hn[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin cVMiV2j8qD0P3CVc315hn[0] <= 16'sb0000000000000000; cVMiV2j8qD0P3CVc315hn[1] <= 16'sb0000000000000000; cVMiV2j8qD0P3CVc315hn[2] <= 16'sb0000000000000000; end else begin cVMiV2j8qD0P3CVc315hn[0] <= a9iZ9svlbzlFdVAGUFPTY[0]; cVMiV2j8qD0P3CVc315hn[1] <= a9iZ9svlbzlFdVAGUFPTY[1]; cVMiV2j8qD0P3CVc315hn[2] <= a9iZ9svlbzlFdVAGUFPTY[2]; end end end assign HeHFnbPrPBgeQHatNQHc0 = cVMiV2j8qD0P3CVc315hn[2]; assign a9iZ9svlbzlFdVAGUFPTY[0] = rFr1ZhZNiURIbPFlZaI4kB; assign a9iZ9svlbzlFdVAGUFPTY[1] = cVMiV2j8qD0P3CVc315hn[0]; assign a9iZ9svlbzlFdVAGUFPTY[2] = cVMiV2j8qD0P3CVc315hn[1]; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : VNPcEW4KZxpAtEz0DCT8vD if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin u2yic2bBqAL2jFtl9bgNqD[0] <= 16'sb0000000000000000; u2yic2bBqAL2jFtl9bgNqD[1] <= 16'sb0000000000000000; u2yic2bBqAL2jFtl9bgNqD[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin u2yic2bBqAL2jFtl9bgNqD[0] <= 16'sb0000000000000000; u2yic2bBqAL2jFtl9bgNqD[1] <= 16'sb0000000000000000; u2yic2bBqAL2jFtl9bgNqD[2] <= 16'sb0000000000000000; end else begin u2yic2bBqAL2jFtl9bgNqD[0] <= rKHf7GW9kd2HwW2mmfwvqC[0]; u2yic2bBqAL2jFtl9bgNqD[1] <= rKHf7GW9kd2HwW2mmfwvqC[1]; u2yic2bBqAL2jFtl9bgNqD[2] <= rKHf7GW9kd2HwW2mmfwvqC[2]; end end end assign gGCeJXlbwaFahBmsH6mMkF = u2yic2bBqAL2jFtl9bgNqD[2]; assign rKHf7GW9kd2HwW2mmfwvqC[0] = gJidztDROiWi1BoJ2KzqKB; assign rKHf7GW9kd2HwW2mmfwvqC[1] = u2yic2bBqAL2jFtl9bgNqD[0]; assign rKHf7GW9kd2HwW2mmfwvqC[2] = u2yic2bBqAL2jFtl9bgNqD[1]; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : t8uWAeIAh3IMbN9UNxoYBKD if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin qM3kFDhftMVWrl1HT1qB4F[0] <= 1'b0; qM3kFDhftMVWrl1HT1qB4F[1] <= 1'b0; qM3kFDhftMVWrl1HT1qB4F[2] <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin qM3kFDhftMVWrl1HT1qB4F[0] <= 1'b0; qM3kFDhftMVWrl1HT1qB4F[1] <= 1'b0; qM3kFDhftMVWrl1HT1qB4F[2] <= 1'b0; end else begin qM3kFDhftMVWrl1HT1qB4F[0] <= eHbdLpdf2r0lFYM9BhuRoB[0]; qM3kFDhftMVWrl1HT1qB4F[1] <= eHbdLpdf2r0lFYM9BhuRoB[1]; qM3kFDhftMVWrl1HT1qB4F[2] <= eHbdLpdf2r0lFYM9BhuRoB[2]; end end end assign l9QVSAqS6jsMaipvGnosLD = qM3kFDhftMVWrl1HT1qB4F[2]; assign eHbdLpdf2r0lFYM9BhuRoB[0] = mm30CTneMiOZJcmmoHkb2D; assign eHbdLpdf2r0lFYM9BhuRoB[1] = qM3kFDhftMVWrl1HT1qB4F[0]; assign eHbdLpdf2r0lFYM9BhuRoB[2] = qM3kFDhftMVWrl1HT1qB4F[1]; cem7BtO0GaQ7W6PGMaiuXF RgLygrKvu632h4sV6s7qoE (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .mm30CTneMiOZJcmmoHkb2D(mm30CTneMiOZJcmmoHkb2D), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .xj58yogg0Lfx8mMLdFuZsE(xj58yogg0Lfx8mMLdFuZsE), .IGbVPdIVOky0HoXMmdGGQH(IGbVPdIVOky0HoXMmdGGQH) ); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : QtzxgwI206U33aXvIkKdwD if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin VzGh5mviLsfsu1Hv3n1l5C <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin VzGh5mviLsfsu1Hv3n1l5C <= 1'b0; end else begin VzGh5mviLsfsu1Hv3n1l5C <= wf5f4XnltnQYt1bEDWEp0F; end end end rjGHdMGdXLgDCNrBAJWf3G mYhLp8wrS9Wo29wMu4jriD (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .FUS5RSCs5VyI8J3rzh0AIE(FUS5RSCs5VyI8J3rzh0AIE), .z8FY0hMnA2CFTR7qvB6dYWC(FUS5RSCs5VyI8J3rzh0AIE), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .g1oJwDFAtNAcPvLahTlMEB(g1oJwDFAtNAcPvLahTlMEB), .wf5f4XnltnQYt1bEDWEp0F(wf5f4XnltnQYt1bEDWEp0F), .Q7D2KKVRLkwEPktPhyCkSD(Q7D2KKVRLkwEPktPhyCkSD) ); htJJjK62gcIcFHavsFtXwE OhCgNBAryg55qaIR7TQ6lD (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .HeHFnbPrPBgeQHatNQHc0(HeHFnbPrPBgeQHatNQHc0), .gGCeJXlbwaFahBmsH6mMkF(gGCeJXlbwaFahBmsH6mMkF), .l9QVSAqS6jsMaipvGnosLD(l9QVSAqS6jsMaipvGnosLD), .g1oJwDFAtNAcPvLahTlMEB(g1oJwDFAtNAcPvLahTlMEB), .VzGh5mviLsfsu1Hv3n1l5C(VzGh5mviLsfsu1Hv3n1l5C), .xj58yogg0Lfx8mMLdFuZsE(xj58yogg0Lfx8mMLdFuZsE), .IGbVPdIVOky0HoXMmdGGQH(IGbVPdIVOky0HoXMmdGGQH), .Q7D2KKVRLkwEPktPhyCkSD(Q7D2KKVRLkwEPktPhyCkSD), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .g1qVkXUxL7Fv5Vq7GJfmGVG(g1qVkXUxL7Fv5Vq7GJfmGVG), .UAWBm55LOUyC0bgEaA5EMC(UAWBm55LOUyC0bgEaA5EMC), .g3JMyJIWtKhpmOxBRsFzIOH(g3JMyJIWtKhpmOxBRsFzIOH), .FUS5RSCs5VyI8J3rzh0AIE(FUS5RSCs5VyI8J3rzh0AIE) ); assign mdal5obekPJm0ao7ZiZ4cF = g1qVkXUxL7Fv5Vq7GJfmGVG; assign j8MMagsoA5t6IysA2ZD3X4F = 1'b1; yzoOoF7555t5sVm5WeZ9lC ZOdIipLNePie2zECiPcAz (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .j8MMagsoA5t6IysA2ZD3X4F(j8MMagsoA5t6IysA2ZD3X4F), .k3VfrgkD6DWITJL9WW5W4D(k3VfrgkD6DWITJL9WW5W4D), .pPn6MVGqBLqJ0xzN2WYfFG(pPn6MVGqBLqJ0xzN2WYfFG), .OUMqBzkN19EDa2VTABMa2E(OUMqBzkN19EDa2VTABMa2E), .qbEnMIxMUsx8pYkF1gFd7D(qbEnMIxMUsx8pYkF1gFd7D), .jNZ4xylBKAANfCL11XNxzB(jNZ4xylBKAANfCL11XNxzB), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .VWSiqDgxQN9a2J7zRy3p4E(aydyoHsGbz0wVGlm34qlsB), .LhqlKpPzANkuN2xC8HYciC(H0BpAwmwCivCDsbLQ5qvCC), .s1N0USypDrc4xyzxc4XEMr(s1N0USypDrc4xyzxc4XEMr), .sZ7bCwrhIAA80IOhzh695(sZ7bCwrhIAA80IOhzh695) ); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : awX33YTQEl2OxkV2HHm04D if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin f69xGE65xXz2LbsT91hgR8G[0] <= 16'sb0000000000000000; f69xGE65xXz2LbsT91hgR8G[1] <= 16'sb0000000000000000; f69xGE65xXz2LbsT91hgR8G[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin f69xGE65xXz2LbsT91hgR8G[0] <= 16'sb0000000000000000; f69xGE65xXz2LbsT91hgR8G[1] <= 16'sb0000000000000000; f69xGE65xXz2LbsT91hgR8G[2] <= 16'sb0000000000000000; end else begin f69xGE65xXz2LbsT91hgR8G[0] <= v4gfbuVl5KUcQzK24qqOvB[0]; f69xGE65xXz2LbsT91hgR8G[1] <= v4gfbuVl5KUcQzK24qqOvB[1]; f69xGE65xXz2LbsT91hgR8G[2] <= v4gfbuVl5KUcQzK24qqOvB[2]; end end end assign DbYwoM2JCYD9mwcRRKmb6G = f69xGE65xXz2LbsT91hgR8G[2]; assign v4gfbuVl5KUcQzK24qqOvB[0] = aydyoHsGbz0wVGlm34qlsB; assign v4gfbuVl5KUcQzK24qqOvB[1] = f69xGE65xXz2LbsT91hgR8G[0]; assign v4gfbuVl5KUcQzK24qqOvB[2] = f69xGE65xXz2LbsT91hgR8G[1]; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : wroVmvZXsLz1H55Ur0PrpB if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin v2G3ZeHqmqPQjfLNmkS0OrG[0] <= 16'sb0000000000000000; v2G3ZeHqmqPQjfLNmkS0OrG[1] <= 16'sb0000000000000000; v2G3ZeHqmqPQjfLNmkS0OrG[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin v2G3ZeHqmqPQjfLNmkS0OrG[0] <= 16'sb0000000000000000; v2G3ZeHqmqPQjfLNmkS0OrG[1] <= 16'sb0000000000000000; v2G3ZeHqmqPQjfLNmkS0OrG[2] <= 16'sb0000000000000000; end else begin v2G3ZeHqmqPQjfLNmkS0OrG[0] <= BrQqlwQZdOtmNiJOrBili[0]; v2G3ZeHqmqPQjfLNmkS0OrG[1] <= BrQqlwQZdOtmNiJOrBili[1]; v2G3ZeHqmqPQjfLNmkS0OrG[2] <= BrQqlwQZdOtmNiJOrBili[2]; end end end assign WbySmFpEqdJe6nrpd6KgG = v2G3ZeHqmqPQjfLNmkS0OrG[2]; assign BrQqlwQZdOtmNiJOrBili[0] = H0BpAwmwCivCDsbLQ5qvCC; assign BrQqlwQZdOtmNiJOrBili[1] = v2G3ZeHqmqPQjfLNmkS0OrG[0]; assign BrQqlwQZdOtmNiJOrBili[2] = v2G3ZeHqmqPQjfLNmkS0OrG[1]; UD63MR6FOodtyKw42f6eiH FYP2YP6G2rKauewwkvNbYC (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .Pq4nKEqqr18aLXK1kX1dfH(Pq4nKEqqr18aLXK1kX1dfH), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .i4y6Td18s9Zr0JbepLQtjC(i4y6Td18s9Zr0JbepLQtjC), .k3FlrGNoOUOhUgHDIDYGouE(k3FlrGNoOUOhUgHDIDYGouE) ); LB48BKt395PB3Xbcuwg3wC w92e99l9cUvs69EuygaxMC (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .DbYwoM2JCYD9mwcRRKmb6G(DbYwoM2JCYD9mwcRRKmb6G), .WbySmFpEqdJe6nrpd6KgG(WbySmFpEqdJe6nrpd6KgG), .pCWATI9lTIGbmXTtLuLAGB(pCWATI9lTIGbmXTtLuLAGB), .yTf5WZbZOLm2uKwJmXk5sG(yTf5WZbZOLm2uKwJmXk5sG), .wGlnEfCkRPxniOjCaZH6XG(wGlnEfCkRPxniOjCaZH6XG), .i4y6Td18s9Zr0JbepLQtjC(i4y6Td18s9Zr0JbepLQtjC), .k3FlrGNoOUOhUgHDIDYGouE(k3FlrGNoOUOhUgHDIDYGouE), .RDvlVEJspE7WkJvNmR8a6C(RDvlVEJspE7WkJvNmR8a6C), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .t30W3eeadZl9O9RnQCafyED(t30W3eeadZl9O9RnQCafyED), .flGpcmOyc38fKmqiV5eQvF(flGpcmOyc38fKmqiV5eQvF) ); TPM8wcrvQfucj4a5DzoryB mrK9eCSSdfMzI9Yt8myOHB (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .t30W3eeadZl9O9RnQCafyED(t30W3eeadZl9O9RnQCafyED), .flGpcmOyc38fKmqiV5eQvF(flGpcmOyc38fKmqiV5eQvF), .DZol1WsbVnSldsei0SiI9E(DZol1WsbVnSldsei0SiI9E), .zqdZMmoxIs9zmnL4kATVuC(zqdZMmoxIs9zmnL4kATVuC), .a8rK4qdEuNCWHLdYbR2f8(a8rK4qdEuNCWHLdYbR2f8), .O6TgnxqnGk692qEmnZQFTC(O6TgnxqnGk692qEmnZQFTC), .XfCDnggI1Y1qaMzSOLL0TD(XfCDnggI1Y1qaMzSOLL0TD), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .CBqrXFTnHQDD2JNQjTxpkH(CBqrXFTnHQDD2JNQjTxpkH), .dYQ3fSOENqw4ZimOQmMMTH(dYQ3fSOENqw4ZimOQmMMTH) ); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : z8NMcVNSFzdoHNpSsC5DBLF if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin k11T3BX1fbEFyiI1W12X7[0] <= 16'sb0000000000000000; k11T3BX1fbEFyiI1W12X7[1] <= 16'sb0000000000000000; k11T3BX1fbEFyiI1W12X7[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin k11T3BX1fbEFyiI1W12X7[0] <= 16'sb0000000000000000; k11T3BX1fbEFyiI1W12X7[1] <= 16'sb0000000000000000; k11T3BX1fbEFyiI1W12X7[2] <= 16'sb0000000000000000; end else begin k11T3BX1fbEFyiI1W12X7[0] <= VpKk1YVVYHSJ6RsO9pshiB[0]; k11T3BX1fbEFyiI1W12X7[1] <= VpKk1YVVYHSJ6RsO9pshiB[1]; k11T3BX1fbEFyiI1W12X7[2] <= VpKk1YVVYHSJ6RsO9pshiB[2]; end end end assign lSTAIQPANZYVi9u1bQJbfC = k11T3BX1fbEFyiI1W12X7[2]; assign VpKk1YVVYHSJ6RsO9pshiB[0] = CBqrXFTnHQDD2JNQjTxpkH; assign VpKk1YVVYHSJ6RsO9pshiB[1] = k11T3BX1fbEFyiI1W12X7[0]; assign VpKk1YVVYHSJ6RsO9pshiB[2] = k11T3BX1fbEFyiI1W12X7[1]; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : j2gHN9roTaQcXLtCUWIL9F if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin RAKTymlGVAtDEhqm1mBWKC[0] <= 16'sb0000000000000000; RAKTymlGVAtDEhqm1mBWKC[1] <= 16'sb0000000000000000; RAKTymlGVAtDEhqm1mBWKC[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin RAKTymlGVAtDEhqm1mBWKC[0] <= 16'sb0000000000000000; RAKTymlGVAtDEhqm1mBWKC[1] <= 16'sb0000000000000000; RAKTymlGVAtDEhqm1mBWKC[2] <= 16'sb0000000000000000; end else begin RAKTymlGVAtDEhqm1mBWKC[0] <= yyMRtRepkZFuqH6zjb0hbC[0]; RAKTymlGVAtDEhqm1mBWKC[1] <= yyMRtRepkZFuqH6zjb0hbC[1]; RAKTymlGVAtDEhqm1mBWKC[2] <= yyMRtRepkZFuqH6zjb0hbC[2]; end end end assign hh7M8p6TyfjHKgE0YxcN3 = RAKTymlGVAtDEhqm1mBWKC[2]; assign yyMRtRepkZFuqH6zjb0hbC[0] = dYQ3fSOENqw4ZimOQmMMTH; assign yyMRtRepkZFuqH6zjb0hbC[1] = RAKTymlGVAtDEhqm1mBWKC[0]; assign yyMRtRepkZFuqH6zjb0hbC[2] = RAKTymlGVAtDEhqm1mBWKC[1]; NdKFdueKdq64dscRK9gG4G k9LBugZcaE827GA1WMmAUmF (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .NMWfejbHi1tIjFkylFWDkC(NMWfejbHi1tIjFkylFWDkC), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .FB6nKajjqrTT1538hBpQ9C(FB6nKajjqrTT1538hBpQ9C), .XcmpMS0nhYnUzTPGBkEmmF(XcmpMS0nhYnUzTPGBkEmmF) ); JRxIvznbGhK1wrungp8WOB rwgHjaAP6nzyxxSYcq7lpF (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .lSTAIQPANZYVi9u1bQJbfC(lSTAIQPANZYVi9u1bQJbfC), .hh7M8p6TyfjHKgE0YxcN3(hh7M8p6TyfjHKgE0YxcN3), .v6PtMRDEb2KzMpzXWCSiwkB(v6PtMRDEb2KzMpzXWCSiwkB), .u6oVvmCf0f079jLPodlV5B(u6oVvmCf0f079jLPodlV5B), .qv4pS1KBm1VYTuOTZHo04F(qv4pS1KBm1VYTuOTZHo04F), .FB6nKajjqrTT1538hBpQ9C(FB6nKajjqrTT1538hBpQ9C), .XcmpMS0nhYnUzTPGBkEmmF(XcmpMS0nhYnUzTPGBkEmmF), .LSv5mOYTPLq5vaIpiVTypC(LSv5mOYTPLq5vaIpiVTypC), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .OAkG388GVoqfAFfrsC3Z3(OAkG388GVoqfAFfrsC3Z3), .DP58bSOk4VSBFH6tnqlVTH(DP58bSOk4VSBFH6tnqlVTH) ); JEVcDj2J0LmsVHIqi6K7z qain7iDZFbUFjqzZeJib6E (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .OAkG388GVoqfAFfrsC3Z3(OAkG388GVoqfAFfrsC3Z3), .DP58bSOk4VSBFH6tnqlVTH(DP58bSOk4VSBFH6tnqlVTH), .Ck459KQ1C8vRbine3lrkt(Ck459KQ1C8vRbine3lrkt), .MCqIdNMOB0Mg1cefHLMjpH(MCqIdNMOB0Mg1cefHLMjpH), .j41GwwL8b9NI9l6ZScQ1PbG(j41GwwL8b9NI9l6ZScQ1PbG), .i8H7HzN3cvjFks6MZ5qaqF(i8H7HzN3cvjFks6MZ5qaqF), .SAcShGLK2YZQrWHGqGVvjD(SAcShGLK2YZQrWHGqGVvjD), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .oEtRmwXRZkMV2JHZdumYM(oEtRmwXRZkMV2JHZdumYM), .ABAJKgUy1j1LH4rwhRtEnG(ABAJKgUy1j1LH4rwhRtEnG) ); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : eVDXDpbSTruDFXBM6ygPaB if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin k9BY0fd7LFxuaZBtnq2NstC[0] <= 16'sb0000000000000000; k9BY0fd7LFxuaZBtnq2NstC[1] <= 16'sb0000000000000000; k9BY0fd7LFxuaZBtnq2NstC[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin k9BY0fd7LFxuaZBtnq2NstC[0] <= 16'sb0000000000000000; k9BY0fd7LFxuaZBtnq2NstC[1] <= 16'sb0000000000000000; k9BY0fd7LFxuaZBtnq2NstC[2] <= 16'sb0000000000000000; end else begin k9BY0fd7LFxuaZBtnq2NstC[0] <= mTZgUkGw3710r8TqEV6XWF[0]; k9BY0fd7LFxuaZBtnq2NstC[1] <= mTZgUkGw3710r8TqEV6XWF[1]; k9BY0fd7LFxuaZBtnq2NstC[2] <= mTZgUkGw3710r8TqEV6XWF[2]; end end end assign PLuy3wDbVIiPXXOVcF7GXC = k9BY0fd7LFxuaZBtnq2NstC[2]; assign mTZgUkGw3710r8TqEV6XWF[0] = oEtRmwXRZkMV2JHZdumYM; assign mTZgUkGw3710r8TqEV6XWF[1] = k9BY0fd7LFxuaZBtnq2NstC[0]; assign mTZgUkGw3710r8TqEV6XWF[2] = k9BY0fd7LFxuaZBtnq2NstC[1]; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : a2bprYW6bhaVvTUhwUfmVQF if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin k8gGlV5iKkuIBPqjsMS5KF[0] <= 16'sb0000000000000000; k8gGlV5iKkuIBPqjsMS5KF[1] <= 16'sb0000000000000000; k8gGlV5iKkuIBPqjsMS5KF[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin k8gGlV5iKkuIBPqjsMS5KF[0] <= 16'sb0000000000000000; k8gGlV5iKkuIBPqjsMS5KF[1] <= 16'sb0000000000000000; k8gGlV5iKkuIBPqjsMS5KF[2] <= 16'sb0000000000000000; end else begin k8gGlV5iKkuIBPqjsMS5KF[0] <= jVudy6rBy3pL4AAajihjvH[0]; k8gGlV5iKkuIBPqjsMS5KF[1] <= jVudy6rBy3pL4AAajihjvH[1]; k8gGlV5iKkuIBPqjsMS5KF[2] <= jVudy6rBy3pL4AAajihjvH[2]; end end end assign wt5uyiFelHvOxXII8I6cTH = k8gGlV5iKkuIBPqjsMS5KF[2]; assign jVudy6rBy3pL4AAajihjvH[0] = ABAJKgUy1j1LH4rwhRtEnG; assign jVudy6rBy3pL4AAajihjvH[1] = k8gGlV5iKkuIBPqjsMS5KF[0]; assign jVudy6rBy3pL4AAajihjvH[2] = k8gGlV5iKkuIBPqjsMS5KF[1]; J3pBieWrBfvDnI3c0xv6sG MwRmE5s9T5vHnHIPrZpBXG (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .mm30CTneMiOZJcmmoHkb2D(mm30CTneMiOZJcmmoHkb2D), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .xj58yogg0Lfx8mMLdFuZsE(gQ8ol00XUcRCyi5uaxpHDB), .IGbVPdIVOky0HoXMmdGGQH(rj0jYY5GSDAuDuCDoIpZ9C) ); I864tK97NgLG3d2RHyF9xG Fd4qoDI1sNmQnnmy3aqxTC (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .HeHFnbPrPBgeQHatNQHc0(PLuy3wDbVIiPXXOVcF7GXC), .gGCeJXlbwaFahBmsH6mMkF(wt5uyiFelHvOxXII8I6cTH), .l9QVSAqS6jsMaipvGnosLD(l9QVSAqS6jsMaipvGnosLD), .g1oJwDFAtNAcPvLahTlMEB(g1oJwDFAtNAcPvLahTlMEB), .VzGh5mviLsfsu1Hv3n1l5C(VzGh5mviLsfsu1Hv3n1l5C), .xj58yogg0Lfx8mMLdFuZsE(gQ8ol00XUcRCyi5uaxpHDB), .IGbVPdIVOky0HoXMmdGGQH(rj0jYY5GSDAuDuCDoIpZ9C), .Q7D2KKVRLkwEPktPhyCkSD(Q7D2KKVRLkwEPktPhyCkSD), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .g1qVkXUxL7Fv5Vq7GJfmGVG(jZwXcJxnQcGGzLJPOScVqE), .UAWBm55LOUyC0bgEaA5EMC(hP5DBuEisrqC9fZ23jziMF) ); assign q4mhS1P9mOTwehAXXNmhxF = jZwXcJxnQcGGzLJPOScVqE; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : RfFhiu7TcZArCuQWZZoVsB if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin x9EdsEkQtjpM4w517iGHzC[0] <= 16'sb0000000000000000; x9EdsEkQtjpM4w517iGHzC[1] <= 16'sb0000000000000000; x9EdsEkQtjpM4w517iGHzC[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin x9EdsEkQtjpM4w517iGHzC[0] <= 16'sb0000000000000000; x9EdsEkQtjpM4w517iGHzC[1] <= 16'sb0000000000000000; x9EdsEkQtjpM4w517iGHzC[2] <= 16'sb0000000000000000; end else begin x9EdsEkQtjpM4w517iGHzC[0] <= tnuZKwedoQlWAtzBo6aIZB[0]; x9EdsEkQtjpM4w517iGHzC[1] <= tnuZKwedoQlWAtzBo6aIZB[1]; x9EdsEkQtjpM4w517iGHzC[2] <= tnuZKwedoQlWAtzBo6aIZB[2]; end end end assign risZnLFYvPBrH1cy6dfHMF = x9EdsEkQtjpM4w517iGHzC[2]; assign tnuZKwedoQlWAtzBo6aIZB[0] = M5AqS9R7rFTkWxwo8io2rH; assign tnuZKwedoQlWAtzBo6aIZB[1] = x9EdsEkQtjpM4w517iGHzC[0]; assign tnuZKwedoQlWAtzBo6aIZB[2] = x9EdsEkQtjpM4w517iGHzC[1]; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : owLoaMKUokO7uUwJJovpJE if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin KmuHj4FutgT59Q7oCiggpD[0] <= 16'sb0000000000000000; KmuHj4FutgT59Q7oCiggpD[1] <= 16'sb0000000000000000; KmuHj4FutgT59Q7oCiggpD[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin KmuHj4FutgT59Q7oCiggpD[0] <= 16'sb0000000000000000; KmuHj4FutgT59Q7oCiggpD[1] <= 16'sb0000000000000000; KmuHj4FutgT59Q7oCiggpD[2] <= 16'sb0000000000000000; end else begin KmuHj4FutgT59Q7oCiggpD[0] <= UFFCUGMTW5jYs8JEV3j3KC[0]; KmuHj4FutgT59Q7oCiggpD[1] <= UFFCUGMTW5jYs8JEV3j3KC[1]; KmuHj4FutgT59Q7oCiggpD[2] <= UFFCUGMTW5jYs8JEV3j3KC[2]; end end end assign y3mUIhc5hpdbI6gB0Klf3MH = KmuHj4FutgT59Q7oCiggpD[2]; assign UFFCUGMTW5jYs8JEV3j3KC[0] = lcJo4MnEaj41ofRAtLkn4D; assign UFFCUGMTW5jYs8JEV3j3KC[1] = KmuHj4FutgT59Q7oCiggpD[0]; assign UFFCUGMTW5jYs8JEV3j3KC[2] = KmuHj4FutgT59Q7oCiggpD[1]; UyxWhYwr5WWgzC84Ncni9D rbo4XnEDAmRflkh99n2moB (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .Pq4nKEqqr18aLXK1kX1dfH(Pq4nKEqqr18aLXK1kX1dfH), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .UlGc2PVtJa9BNobxUHDxSG(UlGc2PVtJa9BNobxUHDxSG), .pdTCH0gTlgy9qR74rtvuBE(pdTCH0gTlgy9qR74rtvuBE) ); wiQ5IhETfzy4iuC7OxoDF ryVcsu5GzuSm41uBLdn2YE (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .risZnLFYvPBrH1cy6dfHMF(risZnLFYvPBrH1cy6dfHMF), .y3mUIhc5hpdbI6gB0Klf3MH(y3mUIhc5hpdbI6gB0Klf3MH), .pCWATI9lTIGbmXTtLuLAGB(pCWATI9lTIGbmXTtLuLAGB), .yTf5WZbZOLm2uKwJmXk5sG(yTf5WZbZOLm2uKwJmXk5sG), .wGlnEfCkRPxniOjCaZH6XG(wGlnEfCkRPxniOjCaZH6XG), .UlGc2PVtJa9BNobxUHDxSG(UlGc2PVtJa9BNobxUHDxSG), .pdTCH0gTlgy9qR74rtvuBE(pdTCH0gTlgy9qR74rtvuBE), .RDvlVEJspE7WkJvNmR8a6C(RDvlVEJspE7WkJvNmR8a6C), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .msLJn85q5aDnigXPSLnA9F(msLJn85q5aDnigXPSLnA9F), .s8tbEDkTdSLkOXc5hVDArH(s8tbEDkTdSLkOXc5hVDArH) ); gOq3QYVANTmyONnNwLvvzB ef4GM1uMXwhosxoRlEdZMF (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .msLJn85q5aDnigXPSLnA9F(msLJn85q5aDnigXPSLnA9F), .s8tbEDkTdSLkOXc5hVDArH(s8tbEDkTdSLkOXc5hVDArH), .DZol1WsbVnSldsei0SiI9E(DZol1WsbVnSldsei0SiI9E), .zqdZMmoxIs9zmnL4kATVuC(zqdZMmoxIs9zmnL4kATVuC), .a8rK4qdEuNCWHLdYbR2f8(a8rK4qdEuNCWHLdYbR2f8), .O6TgnxqnGk692qEmnZQFTC(O6TgnxqnGk692qEmnZQFTC), .XfCDnggI1Y1qaMzSOLL0TD(XfCDnggI1Y1qaMzSOLL0TD), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .ACHpp43jQbQJO4HdGlLQ0B(ACHpp43jQbQJO4HdGlLQ0B), .BJNXQzaMpa7r8LYTHlOrBD(BJNXQzaMpa7r8LYTHlOrBD) ); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : YKhHebQtfFPtGJB8AN9NfC if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin appAG8sqUT59wY8ObKEssF[0] <= 16'sb0000000000000000; appAG8sqUT59wY8ObKEssF[1] <= 16'sb0000000000000000; appAG8sqUT59wY8ObKEssF[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin appAG8sqUT59wY8ObKEssF[0] <= 16'sb0000000000000000; appAG8sqUT59wY8ObKEssF[1] <= 16'sb0000000000000000; appAG8sqUT59wY8ObKEssF[2] <= 16'sb0000000000000000; end else begin appAG8sqUT59wY8ObKEssF[0] <= d21AAbScpxqwLWzuGxj8ajB[0]; appAG8sqUT59wY8ObKEssF[1] <= d21AAbScpxqwLWzuGxj8ajB[1]; appAG8sqUT59wY8ObKEssF[2] <= d21AAbScpxqwLWzuGxj8ajB[2]; end end end assign BXAaMHpKzPpYZGFRqoevNE = appAG8sqUT59wY8ObKEssF[2]; assign d21AAbScpxqwLWzuGxj8ajB[0] = ACHpp43jQbQJO4HdGlLQ0B; assign d21AAbScpxqwLWzuGxj8ajB[1] = appAG8sqUT59wY8ObKEssF[0]; assign d21AAbScpxqwLWzuGxj8ajB[2] = appAG8sqUT59wY8ObKEssF[1]; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : R02gF8dBxGuXtqNBiytOBD if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin pISZVQJtPY1M87J4LAx1MB[0] <= 16'sb0000000000000000; pISZVQJtPY1M87J4LAx1MB[1] <= 16'sb0000000000000000; pISZVQJtPY1M87J4LAx1MB[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin pISZVQJtPY1M87J4LAx1MB[0] <= 16'sb0000000000000000; pISZVQJtPY1M87J4LAx1MB[1] <= 16'sb0000000000000000; pISZVQJtPY1M87J4LAx1MB[2] <= 16'sb0000000000000000; end else begin pISZVQJtPY1M87J4LAx1MB[0] <= EwyTeOtw0Znxv6WUZIsKtH[0]; pISZVQJtPY1M87J4LAx1MB[1] <= EwyTeOtw0Znxv6WUZIsKtH[1]; pISZVQJtPY1M87J4LAx1MB[2] <= EwyTeOtw0Znxv6WUZIsKtH[2]; end end end assign czP63K90EaJdtsY9EHZ30D = pISZVQJtPY1M87J4LAx1MB[2]; assign EwyTeOtw0Znxv6WUZIsKtH[0] = BJNXQzaMpa7r8LYTHlOrBD; assign EwyTeOtw0Znxv6WUZIsKtH[1] = pISZVQJtPY1M87J4LAx1MB[0]; assign EwyTeOtw0Znxv6WUZIsKtH[2] = pISZVQJtPY1M87J4LAx1MB[1]; b3kfX7EdyW6iQU4vGYhPbCG rq8qvMxzcI3hsMYdni7iCG (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .NMWfejbHi1tIjFkylFWDkC(NMWfejbHi1tIjFkylFWDkC), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .mxtJaiWQH83FcZ66WqnMiH(mxtJaiWQH83FcZ66WqnMiH), .MtlWbaE0z2xTCIy368PlWF(MtlWbaE0z2xTCIy368PlWF) ); l9MJ6AwAxJzPDBhrXOVFEiF NueGwXUbsNsksA8LXNYmz (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .BXAaMHpKzPpYZGFRqoevNE(BXAaMHpKzPpYZGFRqoevNE), .czP63K90EaJdtsY9EHZ30D(czP63K90EaJdtsY9EHZ30D), .v6PtMRDEb2KzMpzXWCSiwkB(v6PtMRDEb2KzMpzXWCSiwkB), .u6oVvmCf0f079jLPodlV5B(u6oVvmCf0f079jLPodlV5B), .qv4pS1KBm1VYTuOTZHo04F(qv4pS1KBm1VYTuOTZHo04F), .mxtJaiWQH83FcZ66WqnMiH(mxtJaiWQH83FcZ66WqnMiH), .MtlWbaE0z2xTCIy368PlWF(MtlWbaE0z2xTCIy368PlWF), .LSv5mOYTPLq5vaIpiVTypC(LSv5mOYTPLq5vaIpiVTypC), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .Sek0doTmbyRuabtHW5JKgH(Sek0doTmbyRuabtHW5JKgH), .h4q2yYljVPy2UhMxEpHXfqG(h4q2yYljVPy2UhMxEpHXfqG) ); XDmQpZazz1Q7PrXWDkbfWF yJxVRtqjhNAc0K7yzwOlqF (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .Sek0doTmbyRuabtHW5JKgH(Sek0doTmbyRuabtHW5JKgH), .h4q2yYljVPy2UhMxEpHXfqG(h4q2yYljVPy2UhMxEpHXfqG), .Ck459KQ1C8vRbine3lrkt(Ck459KQ1C8vRbine3lrkt), .MCqIdNMOB0Mg1cefHLMjpH(MCqIdNMOB0Mg1cefHLMjpH), .j41GwwL8b9NI9l6ZScQ1PbG(j41GwwL8b9NI9l6ZScQ1PbG), .i8H7HzN3cvjFks6MZ5qaqF(i8H7HzN3cvjFks6MZ5qaqF), .SAcShGLK2YZQrWHGqGVvjD(SAcShGLK2YZQrWHGqGVvjD), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .Ni5CWVNOepdNWeLhPbktyC(Ni5CWVNOepdNWeLhPbktyC), .oC9IZ8suhbNZiMMpUwYFZE(oC9IZ8suhbNZiMMpUwYFZE) ); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : Fxt9eCqtG0jUXmLi6jZUvE if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin ufyCKBsm7ZcDMoHa9lVT8B[0] <= 16'sb0000000000000000; ufyCKBsm7ZcDMoHa9lVT8B[1] <= 16'sb0000000000000000; ufyCKBsm7ZcDMoHa9lVT8B[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin ufyCKBsm7ZcDMoHa9lVT8B[0] <= 16'sb0000000000000000; ufyCKBsm7ZcDMoHa9lVT8B[1] <= 16'sb0000000000000000; ufyCKBsm7ZcDMoHa9lVT8B[2] <= 16'sb0000000000000000; end else begin ufyCKBsm7ZcDMoHa9lVT8B[0] <= lc0FzXjU6ruJOOuwpT5PQ[0]; ufyCKBsm7ZcDMoHa9lVT8B[1] <= lc0FzXjU6ruJOOuwpT5PQ[1]; ufyCKBsm7ZcDMoHa9lVT8B[2] <= lc0FzXjU6ruJOOuwpT5PQ[2]; end end end assign z6SwcDGEsoURdwbnSfOpHB = ufyCKBsm7ZcDMoHa9lVT8B[2]; assign lc0FzXjU6ruJOOuwpT5PQ[0] = Ni5CWVNOepdNWeLhPbktyC; assign lc0FzXjU6ruJOOuwpT5PQ[1] = ufyCKBsm7ZcDMoHa9lVT8B[0]; assign lc0FzXjU6ruJOOuwpT5PQ[2] = ufyCKBsm7ZcDMoHa9lVT8B[1]; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : iRHyolisTvsKLxVejMexAB if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin f6n0j0rIhtlF1cK7ntOhdG[0] <= 16'sb0000000000000000; f6n0j0rIhtlF1cK7ntOhdG[1] <= 16'sb0000000000000000; f6n0j0rIhtlF1cK7ntOhdG[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin f6n0j0rIhtlF1cK7ntOhdG[0] <= 16'sb0000000000000000; f6n0j0rIhtlF1cK7ntOhdG[1] <= 16'sb0000000000000000; f6n0j0rIhtlF1cK7ntOhdG[2] <= 16'sb0000000000000000; end else begin f6n0j0rIhtlF1cK7ntOhdG[0] <= f8PGb7nqRvYgidEKAnbVYCF[0]; f6n0j0rIhtlF1cK7ntOhdG[1] <= f8PGb7nqRvYgidEKAnbVYCF[1]; f6n0j0rIhtlF1cK7ntOhdG[2] <= f8PGb7nqRvYgidEKAnbVYCF[2]; end end end assign pGKHaOZvJloUuxOXANTYZE = f6n0j0rIhtlF1cK7ntOhdG[2]; assign f8PGb7nqRvYgidEKAnbVYCF[0] = oC9IZ8suhbNZiMMpUwYFZE; assign f8PGb7nqRvYgidEKAnbVYCF[1] = f6n0j0rIhtlF1cK7ntOhdG[0]; assign f8PGb7nqRvYgidEKAnbVYCF[2] = f6n0j0rIhtlF1cK7ntOhdG[1]; B4aNKopc1IycejU6cc0njB bQVBAnxXJylfCrtgM5vSPE (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .mm30CTneMiOZJcmmoHkb2D(mm30CTneMiOZJcmmoHkb2D), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .xj58yogg0Lfx8mMLdFuZsE(feyfHDrrhsk9bdeB57O2c), .IGbVPdIVOky0HoXMmdGGQH(r2IKtvrSH76nVotfMIojNdD) ); nma7TM3OXSEWWsbewMlcHG m3c8ml2wLBYxENxWE5xJzkC (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .HeHFnbPrPBgeQHatNQHc0(z6SwcDGEsoURdwbnSfOpHB), .gGCeJXlbwaFahBmsH6mMkF(pGKHaOZvJloUuxOXANTYZE), .l9QVSAqS6jsMaipvGnosLD(l9QVSAqS6jsMaipvGnosLD), .g1oJwDFAtNAcPvLahTlMEB(g1oJwDFAtNAcPvLahTlMEB), .VzGh5mviLsfsu1Hv3n1l5C(VzGh5mviLsfsu1Hv3n1l5C), .xj58yogg0Lfx8mMLdFuZsE(feyfHDrrhsk9bdeB57O2c), .IGbVPdIVOky0HoXMmdGGQH(r2IKtvrSH76nVotfMIojNdD), .Q7D2KKVRLkwEPktPhyCkSD(Q7D2KKVRLkwEPktPhyCkSD), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .g1qVkXUxL7Fv5Vq7GJfmGVG(SmUoeWULdUSlbsjccscXpG), .UAWBm55LOUyC0bgEaA5EMC(qrJeNpaPfOy0pMCu40c1ME) ); assign vyWRmDyKy2RVVIdRBtzV5F = SmUoeWULdUSlbsjccscXpG; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : e6AZe9KIcZJURxtpakQhtqG if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin hDe4KgCGLUE2lc3mBRHUGE[0] <= 16'sb0000000000000000; hDe4KgCGLUE2lc3mBRHUGE[1] <= 16'sb0000000000000000; hDe4KgCGLUE2lc3mBRHUGE[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin hDe4KgCGLUE2lc3mBRHUGE[0] <= 16'sb0000000000000000; hDe4KgCGLUE2lc3mBRHUGE[1] <= 16'sb0000000000000000; hDe4KgCGLUE2lc3mBRHUGE[2] <= 16'sb0000000000000000; end else begin hDe4KgCGLUE2lc3mBRHUGE[0] <= ZvqDLDMtFPbHpUtzihpbXF[0]; hDe4KgCGLUE2lc3mBRHUGE[1] <= ZvqDLDMtFPbHpUtzihpbXF[1]; hDe4KgCGLUE2lc3mBRHUGE[2] <= ZvqDLDMtFPbHpUtzihpbXF[2]; end end end assign EiKTmNA9gqnqt6QU2ytsGF = hDe4KgCGLUE2lc3mBRHUGE[2]; assign ZvqDLDMtFPbHpUtzihpbXF[0] = s1N0USypDrc4xyzxc4XEMr; assign ZvqDLDMtFPbHpUtzihpbXF[1] = hDe4KgCGLUE2lc3mBRHUGE[0]; assign ZvqDLDMtFPbHpUtzihpbXF[2] = hDe4KgCGLUE2lc3mBRHUGE[1]; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : y8LVueovJyghRSuIm8a5QH if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin I3TwcvTY4hEZBUKyNKGQYH[0] <= 16'sb0000000000000000; I3TwcvTY4hEZBUKyNKGQYH[1] <= 16'sb0000000000000000; I3TwcvTY4hEZBUKyNKGQYH[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin I3TwcvTY4hEZBUKyNKGQYH[0] <= 16'sb0000000000000000; I3TwcvTY4hEZBUKyNKGQYH[1] <= 16'sb0000000000000000; I3TwcvTY4hEZBUKyNKGQYH[2] <= 16'sb0000000000000000; end else begin I3TwcvTY4hEZBUKyNKGQYH[0] <= ltutKZEJ3uAsYBtveZfxN[0]; I3TwcvTY4hEZBUKyNKGQYH[1] <= ltutKZEJ3uAsYBtveZfxN[1]; I3TwcvTY4hEZBUKyNKGQYH[2] <= ltutKZEJ3uAsYBtveZfxN[2]; end end end assign i0padod73DFvzROjA4fS2o = I3TwcvTY4hEZBUKyNKGQYH[2]; assign ltutKZEJ3uAsYBtveZfxN[0] = sZ7bCwrhIAA80IOhzh695; assign ltutKZEJ3uAsYBtveZfxN[1] = I3TwcvTY4hEZBUKyNKGQYH[0]; assign ltutKZEJ3uAsYBtveZfxN[2] = I3TwcvTY4hEZBUKyNKGQYH[1]; q2kRA8XOHHRNcp89kCO6bC I2TBaFHPkLkB0woW45YSD (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .Pq4nKEqqr18aLXK1kX1dfH(Pq4nKEqqr18aLXK1kX1dfH), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .mvb8xVo6CcFPFyQu3ctDE(mvb8xVo6CcFPFyQu3ctDE), .gC05dypmmuscVux3EfDHCD(gC05dypmmuscVux3EfDHCD) ); zkst6F43f7ijCyz44loHhB t9g2Y8fM4yk65azUUSe1E3F (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .EiKTmNA9gqnqt6QU2ytsGF(EiKTmNA9gqnqt6QU2ytsGF), .i0padod73DFvzROjA4fS2o(i0padod73DFvzROjA4fS2o), .pCWATI9lTIGbmXTtLuLAGB(pCWATI9lTIGbmXTtLuLAGB), .yTf5WZbZOLm2uKwJmXk5sG(yTf5WZbZOLm2uKwJmXk5sG), .wGlnEfCkRPxniOjCaZH6XG(wGlnEfCkRPxniOjCaZH6XG), .mvb8xVo6CcFPFyQu3ctDE(mvb8xVo6CcFPFyQu3ctDE), .gC05dypmmuscVux3EfDHCD(gC05dypmmuscVux3EfDHCD), .RDvlVEJspE7WkJvNmR8a6C(RDvlVEJspE7WkJvNmR8a6C), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .DxKKPTJNNNGcVbnDyBefdC(DxKKPTJNNNGcVbnDyBefdC), .z5IVnN9scVD1jMboeUZaZG(z5IVnN9scVD1jMboeUZaZG) ); bXwzfDHB1o41csk9RIaLuD bY2yqF5WO84iCOvXu7u5gH (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .DxKKPTJNNNGcVbnDyBefdC(DxKKPTJNNNGcVbnDyBefdC), .z5IVnN9scVD1jMboeUZaZG(z5IVnN9scVD1jMboeUZaZG), .DZol1WsbVnSldsei0SiI9E(DZol1WsbVnSldsei0SiI9E), .zqdZMmoxIs9zmnL4kATVuC(zqdZMmoxIs9zmnL4kATVuC), .a8rK4qdEuNCWHLdYbR2f8(a8rK4qdEuNCWHLdYbR2f8), .O6TgnxqnGk692qEmnZQFTC(O6TgnxqnGk692qEmnZQFTC), .XfCDnggI1Y1qaMzSOLL0TD(XfCDnggI1Y1qaMzSOLL0TD), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .y2F62Qir2uvIcDNjqoCgbPG(y2F62Qir2uvIcDNjqoCgbPG), .eJSHu1mAvW9BzbMy0ufWWD(eJSHu1mAvW9BzbMy0ufWWD) ); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : Yera4SjAVuKG7TjeL0xum if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin h41dWYc0X3ZAsDk44FMtsTD[0] <= 16'sb0000000000000000; h41dWYc0X3ZAsDk44FMtsTD[1] <= 16'sb0000000000000000; h41dWYc0X3ZAsDk44FMtsTD[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin h41dWYc0X3ZAsDk44FMtsTD[0] <= 16'sb0000000000000000; h41dWYc0X3ZAsDk44FMtsTD[1] <= 16'sb0000000000000000; h41dWYc0X3ZAsDk44FMtsTD[2] <= 16'sb0000000000000000; end else begin h41dWYc0X3ZAsDk44FMtsTD[0] <= kZIaatjtNR5S1owTPfmSI[0]; h41dWYc0X3ZAsDk44FMtsTD[1] <= kZIaatjtNR5S1owTPfmSI[1]; h41dWYc0X3ZAsDk44FMtsTD[2] <= kZIaatjtNR5S1owTPfmSI[2]; end end end assign SNl44VPeKmo2uIh5zCljYE = h41dWYc0X3ZAsDk44FMtsTD[2]; assign kZIaatjtNR5S1owTPfmSI[0] = y2F62Qir2uvIcDNjqoCgbPG; assign kZIaatjtNR5S1owTPfmSI[1] = h41dWYc0X3ZAsDk44FMtsTD[0]; assign kZIaatjtNR5S1owTPfmSI[2] = h41dWYc0X3ZAsDk44FMtsTD[1]; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : MplkH2AOPP4uw14V7wrk3B if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin UbhppxZFtuRiGSMYxgMT2F[0] <= 16'sb0000000000000000; UbhppxZFtuRiGSMYxgMT2F[1] <= 16'sb0000000000000000; UbhppxZFtuRiGSMYxgMT2F[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin UbhppxZFtuRiGSMYxgMT2F[0] <= 16'sb0000000000000000; UbhppxZFtuRiGSMYxgMT2F[1] <= 16'sb0000000000000000; UbhppxZFtuRiGSMYxgMT2F[2] <= 16'sb0000000000000000; end else begin UbhppxZFtuRiGSMYxgMT2F[0] <= rk6XtqxIQmYnoKIvpO9PNH[0]; UbhppxZFtuRiGSMYxgMT2F[1] <= rk6XtqxIQmYnoKIvpO9PNH[1]; UbhppxZFtuRiGSMYxgMT2F[2] <= rk6XtqxIQmYnoKIvpO9PNH[2]; end end end assign AXkTVaeFKW3Cvod76gwXK = UbhppxZFtuRiGSMYxgMT2F[2]; assign rk6XtqxIQmYnoKIvpO9PNH[0] = eJSHu1mAvW9BzbMy0ufWWD; assign rk6XtqxIQmYnoKIvpO9PNH[1] = UbhppxZFtuRiGSMYxgMT2F[0]; assign rk6XtqxIQmYnoKIvpO9PNH[2] = UbhppxZFtuRiGSMYxgMT2F[1]; AMV8VvUfHFpyXwL05KB5KG jZAgC07ng8reotvX6puRbG (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .NMWfejbHi1tIjFkylFWDkC(NMWfejbHi1tIjFkylFWDkC), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .PV2GPYF9MTfm6A3VIE3yL(PV2GPYF9MTfm6A3VIE3yL), .VMMfdu9AIUdQe4XcwZLbSC(VMMfdu9AIUdQe4XcwZLbSC) ); yJ9pGr1LKI77BCyDbnt2UC x9yUjJ4dQaL4JCZ6bTAoBB (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .SNl44VPeKmo2uIh5zCljYE(SNl44VPeKmo2uIh5zCljYE), .AXkTVaeFKW3Cvod76gwXK(AXkTVaeFKW3Cvod76gwXK), .v6PtMRDEb2KzMpzXWCSiwkB(v6PtMRDEb2KzMpzXWCSiwkB), .u6oVvmCf0f079jLPodlV5B(u6oVvmCf0f079jLPodlV5B), .qv4pS1KBm1VYTuOTZHo04F(qv4pS1KBm1VYTuOTZHo04F), .PV2GPYF9MTfm6A3VIE3yL(PV2GPYF9MTfm6A3VIE3yL), .VMMfdu9AIUdQe4XcwZLbSC(VMMfdu9AIUdQe4XcwZLbSC), .LSv5mOYTPLq5vaIpiVTypC(LSv5mOYTPLq5vaIpiVTypC), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .BSA6wYLjrd40iGAxWAWPUG(BSA6wYLjrd40iGAxWAWPUG), .mVsThSJWeEPGLaZQZJ476C(mVsThSJWeEPGLaZQZJ476C) ); rjG8zPr4pPV2nTcp1wQ6sE frmFPr2Hgpf7JABWVreFmH (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .BSA6wYLjrd40iGAxWAWPUG(BSA6wYLjrd40iGAxWAWPUG), .mVsThSJWeEPGLaZQZJ476C(mVsThSJWeEPGLaZQZJ476C), .Ck459KQ1C8vRbine3lrkt(Ck459KQ1C8vRbine3lrkt), .MCqIdNMOB0Mg1cefHLMjpH(MCqIdNMOB0Mg1cefHLMjpH), .j41GwwL8b9NI9l6ZScQ1PbG(j41GwwL8b9NI9l6ZScQ1PbG), .i8H7HzN3cvjFks6MZ5qaqF(i8H7HzN3cvjFks6MZ5qaqF), .SAcShGLK2YZQrWHGqGVvjD(SAcShGLK2YZQrWHGqGVvjD), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .Qjop49qrCNJ2RVI1tmxWK(Qjop49qrCNJ2RVI1tmxWK), .qtlf3VUxsnDXMsfKMVqqRD(qtlf3VUxsnDXMsfKMVqqRD) ); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : QkTsAMX2ysQgjvkiAUs2oC if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin TGSVeodh4aSh5YMUFsJBpF[0] <= 16'sb0000000000000000; TGSVeodh4aSh5YMUFsJBpF[1] <= 16'sb0000000000000000; TGSVeodh4aSh5YMUFsJBpF[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin TGSVeodh4aSh5YMUFsJBpF[0] <= 16'sb0000000000000000; TGSVeodh4aSh5YMUFsJBpF[1] <= 16'sb0000000000000000; TGSVeodh4aSh5YMUFsJBpF[2] <= 16'sb0000000000000000; end else begin TGSVeodh4aSh5YMUFsJBpF[0] <= pKwMCjbBuwX4wlYrJtZeqH[0]; TGSVeodh4aSh5YMUFsJBpF[1] <= pKwMCjbBuwX4wlYrJtZeqH[1]; TGSVeodh4aSh5YMUFsJBpF[2] <= pKwMCjbBuwX4wlYrJtZeqH[2]; end end end assign T6wR1FRvpbz8HFANbQ6odH = TGSVeodh4aSh5YMUFsJBpF[2]; assign pKwMCjbBuwX4wlYrJtZeqH[0] = Qjop49qrCNJ2RVI1tmxWK; assign pKwMCjbBuwX4wlYrJtZeqH[1] = TGSVeodh4aSh5YMUFsJBpF[0]; assign pKwMCjbBuwX4wlYrJtZeqH[2] = TGSVeodh4aSh5YMUFsJBpF[1]; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : EUqbtBsMjpkspgfBj9UDCG if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin t1XxIWfdmuGYgMJ14AA5aoF[0] <= 16'sb0000000000000000; t1XxIWfdmuGYgMJ14AA5aoF[1] <= 16'sb0000000000000000; t1XxIWfdmuGYgMJ14AA5aoF[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin t1XxIWfdmuGYgMJ14AA5aoF[0] <= 16'sb0000000000000000; t1XxIWfdmuGYgMJ14AA5aoF[1] <= 16'sb0000000000000000; t1XxIWfdmuGYgMJ14AA5aoF[2] <= 16'sb0000000000000000; end else begin t1XxIWfdmuGYgMJ14AA5aoF[0] <= Ed8ZUSDNSkOaxlQSyerJMG[0]; t1XxIWfdmuGYgMJ14AA5aoF[1] <= Ed8ZUSDNSkOaxlQSyerJMG[1]; t1XxIWfdmuGYgMJ14AA5aoF[2] <= Ed8ZUSDNSkOaxlQSyerJMG[2]; end end end assign c88iPPDCYH3uMXl21XZoi8D = t1XxIWfdmuGYgMJ14AA5aoF[2]; assign Ed8ZUSDNSkOaxlQSyerJMG[0] = qtlf3VUxsnDXMsfKMVqqRD; assign Ed8ZUSDNSkOaxlQSyerJMG[1] = t1XxIWfdmuGYgMJ14AA5aoF[0]; assign Ed8ZUSDNSkOaxlQSyerJMG[2] = t1XxIWfdmuGYgMJ14AA5aoF[1]; x0QNWtVHJg3u2GVrxFhqr7C F90JVXWaKZWqArerfGE6dF (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .mm30CTneMiOZJcmmoHkb2D(mm30CTneMiOZJcmmoHkb2D), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .xj58yogg0Lfx8mMLdFuZsE(RRE1h6KsUsyxLABwNoPOPB), .IGbVPdIVOky0HoXMmdGGQH(vM9w9urjKvIy07zqFkMIPF) ); h6yzizqXIBvb7BHvowGhhgB Zej2MHUlV16aYtNg9H5IsC (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .HeHFnbPrPBgeQHatNQHc0(T6wR1FRvpbz8HFANbQ6odH), .gGCeJXlbwaFahBmsH6mMkF(c88iPPDCYH3uMXl21XZoi8D), .l9QVSAqS6jsMaipvGnosLD(l9QVSAqS6jsMaipvGnosLD), .g1oJwDFAtNAcPvLahTlMEB(g1oJwDFAtNAcPvLahTlMEB), .VzGh5mviLsfsu1Hv3n1l5C(VzGh5mviLsfsu1Hv3n1l5C), .xj58yogg0Lfx8mMLdFuZsE(RRE1h6KsUsyxLABwNoPOPB), .IGbVPdIVOky0HoXMmdGGQH(vM9w9urjKvIy07zqFkMIPF), .Q7D2KKVRLkwEPktPhyCkSD(Q7D2KKVRLkwEPktPhyCkSD), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .g1qVkXUxL7Fv5Vq7GJfmGVG(tZCSNlfV8pGx0wl9RXazqC), .UAWBm55LOUyC0bgEaA5EMC(vuJEKfnV5iqg56DSJMMzfH) ); assign SRoFC9yIIwEIUwYpoyy0QF = tZCSNlfV8pGx0wl9RXazqC; assign wpHiLzmis5ns3l38MddOzE = UAWBm55LOUyC0bgEaA5EMC; assign j963sPBld8mpm71sqcvb8WF = hP5DBuEisrqC9fZ23jziMF; assign Ic4vfYy6jnxaw8uXI98INH = qrJeNpaPfOy0pMCu40c1ME; assign x2KkW4HKTQgVBmVskDu4RD = vuJEKfnV5iqg56DSJMMzfH; assign g1D8wSsV4Ksuy5G0qxKYMs = g3JMyJIWtKhpmOxBRsFzIOH; endmodule