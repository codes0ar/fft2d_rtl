`timescale 1 ns / 1 ns module am04sFwquwsZE10aTKfoWG (v04pHKxyc2sPW047bbyUgE, JAMOfrNHxGSYDF0urqkLN, IPh1M0O3x0ioGlon72MROG, Mt05SNCQbo0cCPNa1yEFyF, xYJCS7zMCKI1yYR3Bx1XrD, AaqUpSvCGAV1YR86nIsLWH, Z7ZDy0EvwvoCh1zahAqvSF, R6zf5iqRNVEGVBO8egq8kF, VWSiqDgxQN9a2J7zRy3p4E, LhqlKpPzANkuN2xC8HYciC, OUMqBzkN19EDa2VTABMa2E, qbEnMIxMUsx8pYkF1gFd7D); input v04pHKxyc2sPW047bbyUgE; input JAMOfrNHxGSYDF0urqkLN; input signed [15:0] IPh1M0O3x0ioGlon72MROG; input signed [15:0] Mt05SNCQbo0cCPNa1yEFyF; input signed [15:0] xYJCS7zMCKI1yYR3Bx1XrD; input signed [15:0] AaqUpSvCGAV1YR86nIsLWH; input Z7ZDy0EvwvoCh1zahAqvSF; input R6zf5iqRNVEGVBO8egq8kF; output signed [15:0] VWSiqDgxQN9a2J7zRy3p4E; output signed [15:0] LhqlKpPzANkuN2xC8HYciC; output signed [15:0] OUMqBzkN19EDa2VTABMa2E; output signed [15:0] qbEnMIxMUsx8pYkF1gFd7D; reg signed [16:0] JuEdAzP84rg2g9z7jUH4CD; reg signed [16:0] w13lDdnHeKbz12RPLclXaYB; reg signed [16:0] G1cI3X0rnsuzwQl9n17YG; reg signed [16:0] GXg6LN8xFsDjdENYEDgKvC; reg c4yitNmVtLmJQVcYGJPLIKF; reg signed [16:0] EwpgnQRNtLL4vjPMlLBwS; reg signed [16:0] wf6CdozoYkNBecSlGbH3aH; reg signed [16:0] EVnidbw743875wavOVIR7C; reg signed [16:0] o238XHbXd6S5MNKr5zezYE; reg u3HkQauhqeq4XUajUjEhKC; reg signed [15:0] aydyoHsGbz0wVGlm34qlsB; reg signed [15:0] H0BpAwmwCivCDsbLQ5qvCC; reg signed [15:0] s1N0USypDrc4xyzxc4XEMr; reg signed [15:0] sZ7bCwrhIAA80IOhzh695; reg ODhxEeLGlzFMjyKZKgHvLB; reg signed [16:0] sePOIYBEAAbt3DPar8jd5F; reg signed [16:0] iR0ShkyVRkHalUKTDnP0tG; reg signed [16:0] j3ureEigNPclVAPr6VwHVbG; reg signed [16:0] PmhJP7JCYGM2OStQXGIHgD; reg signed [16:0] TqfF3Zgxtm2cKWvwqij3m; reg signed [16:0] xijHKILnnZ8AgezrLRQvfF; reg signed [16:0] LoYaOvLnEQPAYlYtjywSTF; reg signed [16:0] Wf2SXd0xW1vBpZ49DhpQPE; reg signed [16:0] q5X9uuOdY7IBIroLr9svCOD; reg signed [16:0] BWK9w55Ml1WM8fecaddoXH; reg signed [16:0] h5B5oTxicZ5M23LhruZny; reg signed [16:0] DZuRxUKTwIbTxoU1h9ItHG; reg signed [16:0] pePHH82YpiwDZXNTNuW0kE; reg signed [16:0] w2JsFHlps9UnWS2sz8ntdrD; reg signed [16:0] Tyt8bZLXYY8su2Ax3b0rDH; reg signed [16:0] FZwXLiG4fwR5D6OFWbauRD; reg signed [16:0] b9TGb0JMaIybP28lLxuqbSD; reg signed [16:0] soGohDPw7ZeleH1CUwdFeD; reg signed [16:0] B8FsciuTU1IBtwPIKxFjdD; reg signed [16:0] V38Q9K9It91xb35KJJQllB; wire J5bxDbhUXfqtoh3x3px8OH; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : cByCCMbEZEcgRtZNjjMl3D if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin JuEdAzP84rg2g9z7jUH4CD <= 17'sb00000000000000000; w13lDdnHeKbz12RPLclXaYB <= 17'sb00000000000000000; G1cI3X0rnsuzwQl9n17YG <= 17'sb00000000000000000; GXg6LN8xFsDjdENYEDgKvC <= 17'sb00000000000000000; c4yitNmVtLmJQVcYGJPLIKF <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin JuEdAzP84rg2g9z7jUH4CD <= 17'sb00000000000000000; w13lDdnHeKbz12RPLclXaYB <= 17'sb00000000000000000; G1cI3X0rnsuzwQl9n17YG <= 17'sb00000000000000000; GXg6LN8xFsDjdENYEDgKvC <= 17'sb00000000000000000; c4yitNmVtLmJQVcYGJPLIKF <= 1'b0; end else begin JuEdAzP84rg2g9z7jUH4CD <= EwpgnQRNtLL4vjPMlLBwS; w13lDdnHeKbz12RPLclXaYB <= wf6CdozoYkNBecSlGbH3aH; G1cI3X0rnsuzwQl9n17YG <= EVnidbw743875wavOVIR7C; GXg6LN8xFsDjdENYEDgKvC <= o238XHbXd6S5MNKr5zezYE; c4yitNmVtLmJQVcYGJPLIKF <= u3HkQauhqeq4XUajUjEhKC; end end end always @(AaqUpSvCGAV1YR86nIsLWH, G1cI3X0rnsuzwQl9n17YG, GXg6LN8xFsDjdENYEDgKvC, IPh1M0O3x0ioGlon72MROG, JuEdAzP84rg2g9z7jUH4CD, Mt05SNCQbo0cCPNa1yEFyF, Z7ZDy0EvwvoCh1zahAqvSF, c4yitNmVtLmJQVcYGJPLIKF, w13lDdnHeKbz12RPLclXaYB, xYJCS7zMCKI1yYR3Bx1XrD) begin pePHH82YpiwDZXNTNuW0kE = 17'sb00000000000000000; w2JsFHlps9UnWS2sz8ntdrD = 17'sb00000000000000000; Tyt8bZLXYY8su2Ax3b0rDH = 17'sb00000000000000000; FZwXLiG4fwR5D6OFWbauRD = 17'sb00000000000000000; b9TGb0JMaIybP28lLxuqbSD = 17'sb00000000000000000; soGohDPw7ZeleH1CUwdFeD = 17'sb00000000000000000; B8FsciuTU1IBtwPIKxFjdD = 17'sb00000000000000000; V38Q9K9It91xb35KJJQllB = 17'sb00000000000000000; EwpgnQRNtLL4vjPMlLBwS = JuEdAzP84rg2g9z7jUH4CD; wf6CdozoYkNBecSlGbH3aH = w13lDdnHeKbz12RPLclXaYB; EVnidbw743875wavOVIR7C = G1cI3X0rnsuzwQl9n17YG; o238XHbXd6S5MNKr5zezYE = GXg6LN8xFsDjdENYEDgKvC; u3HkQauhqeq4XUajUjEhKC = Z7ZDy0EvwvoCh1zahAqvSF; if (Z7ZDy0EvwvoCh1zahAqvSF) begin pePHH82YpiwDZXNTNuW0kE = {IPh1M0O3x0ioGlon72MROG[15], IPh1M0O3x0ioGlon72MROG}; w2JsFHlps9UnWS2sz8ntdrD = {xYJCS7zMCKI1yYR3Bx1XrD[15], xYJCS7zMCKI1yYR3Bx1XrD}; EwpgnQRNtLL4vjPMlLBwS = pePHH82YpiwDZXNTNuW0kE + w2JsFHlps9UnWS2sz8ntdrD; Tyt8bZLXYY8su2Ax3b0rDH = {IPh1M0O3x0ioGlon72MROG[15], IPh1M0O3x0ioGlon72MROG}; FZwXLiG4fwR5D6OFWbauRD = {xYJCS7zMCKI1yYR3Bx1XrD[15], xYJCS7zMCKI1yYR3Bx1XrD}; EVnidbw743875wavOVIR7C = Tyt8bZLXYY8su2Ax3b0rDH - FZwXLiG4fwR5D6OFWbauRD; b9TGb0JMaIybP28lLxuqbSD = {Mt05SNCQbo0cCPNa1yEFyF[15], Mt05SNCQbo0cCPNa1yEFyF}; soGohDPw7ZeleH1CUwdFeD = {AaqUpSvCGAV1YR86nIsLWH[15], AaqUpSvCGAV1YR86nIsLWH}; wf6CdozoYkNBecSlGbH3aH = b9TGb0JMaIybP28lLxuqbSD + soGohDPw7ZeleH1CUwdFeD; B8FsciuTU1IBtwPIKxFjdD = {Mt05SNCQbo0cCPNa1yEFyF[15], Mt05SNCQbo0cCPNa1yEFyF}; V38Q9K9It91xb35KJJQllB = {AaqUpSvCGAV1YR86nIsLWH[15], AaqUpSvCGAV1YR86nIsLWH}; o238XHbXd6S5MNKr5zezYE = B8FsciuTU1IBtwPIKxFjdD - V38Q9K9It91xb35KJJQllB; end sePOIYBEAAbt3DPar8jd5F = ({JuEdAzP84rg2g9z7jUH4CD[16], JuEdAzP84rg2g9z7jUH4CD[16:1]}) + $signed({1'b0, JuEdAzP84rg2g9z7jUH4CD[0]}); iR0ShkyVRkHalUKTDnP0tG = sePOIYBEAAbt3DPar8jd5F >>> 8'd1; j3ureEigNPclVAPr6VwHVbG = {iR0ShkyVRkHalUKTDnP0tG[15:0], 1'b0}; aydyoHsGbz0wVGlm34qlsB = j3ureEigNPclVAPr6VwHVbG[15:0]; PmhJP7JCYGM2OStQXGIHgD = ({w13lDdnHeKbz12RPLclXaYB[16], w13lDdnHeKbz12RPLclXaYB[16:1]}) + $signed({1'b0, w13lDdnHeKbz12RPLclXaYB[0]}); TqfF3Zgxtm2cKWvwqij3m = PmhJP7JCYGM2OStQXGIHgD >>> 8'd1; xijHKILnnZ8AgezrLRQvfF = {TqfF3Zgxtm2cKWvwqij3m[15:0], 1'b0}; H0BpAwmwCivCDsbLQ5qvCC = xijHKILnnZ8AgezrLRQvfF[15:0]; LoYaOvLnEQPAYlYtjywSTF = ({G1cI3X0rnsuzwQl9n17YG[16], G1cI3X0rnsuzwQl9n17YG[16:1]}) + $signed({1'b0, G1cI3X0rnsuzwQl9n17YG[0]}); Wf2SXd0xW1vBpZ49DhpQPE = LoYaOvLnEQPAYlYtjywSTF >>> 8'd1; q5X9uuOdY7IBIroLr9svCOD = {Wf2SXd0xW1vBpZ49DhpQPE[15:0], 1'b0}; s1N0USypDrc4xyzxc4XEMr = q5X9uuOdY7IBIroLr9svCOD[15:0]; BWK9w55Ml1WM8fecaddoXH = ({GXg6LN8xFsDjdENYEDgKvC[16], GXg6LN8xFsDjdENYEDgKvC[16:1]}) + $signed({1'b0, GXg6LN8xFsDjdENYEDgKvC[0]}); h5B5oTxicZ5M23LhruZny = BWK9w55Ml1WM8fecaddoXH >>> 8'd1; DZuRxUKTwIbTxoU1h9ItHG = {h5B5oTxicZ5M23LhruZny[15:0], 1'b0}; sZ7bCwrhIAA80IOhzh695 = DZuRxUKTwIbTxoU1h9ItHG[15:0]; ODhxEeLGlzFMjyKZKgHvLB = c4yitNmVtLmJQVcYGJPLIKF; end assign VWSiqDgxQN9a2J7zRy3p4E = aydyoHsGbz0wVGlm34qlsB; assign LhqlKpPzANkuN2xC8HYciC = H0BpAwmwCivCDsbLQ5qvCC; assign OUMqBzkN19EDa2VTABMa2E = s1N0USypDrc4xyzxc4XEMr; assign qbEnMIxMUsx8pYkF1gFd7D = sZ7bCwrhIAA80IOhzh695; endmodule