`timescale 1 ns / 1 ns module QNagGs9mRrlwXRNR72KVyF (v04pHKxyc2sPW047bbyUgE, JAMOfrNHxGSYDF0urqkLN, Ck459KQ1C8vRbine3lrkt, DCqZJgzh8RI4wgf1TYRoc, R6zf5iqRNVEGVBO8egq8kF, MCqIdNMOB0Mg1cefHLMjpH, j41GwwL8b9NI9l6ZScQ1PbG, i8H7HzN3cvjFks6MZ5qaqF, SAcShGLK2YZQrWHGqGVvjD); input v04pHKxyc2sPW047bbyUgE; input JAMOfrNHxGSYDF0urqkLN; input Ck459KQ1C8vRbine3lrkt; input DCqZJgzh8RI4wgf1TYRoc; input R6zf5iqRNVEGVBO8egq8kF; output [2:0] MCqIdNMOB0Mg1cefHLMjpH; output j41GwwL8b9NI9l6ZScQ1PbG; output i8H7HzN3cvjFks6MZ5qaqF; output SAcShGLK2YZQrWHGqGVvjD; reg [2:0] JomiEQo6ylRrlhLJPFsQTG; reg [1:0] X7FJ0jgk6hqdMN8BingGvE; reg [1:0] WXS42gmgDxS46057b3AGD; reg [2:0] GP01IUV0xObQQCSdqL463C; reg pDYTWTp6fyrEdA1XnDiP6E; reg [1:0] mb13NdjIe7rpJDLNih8AaE; reg Xf88wK4mkniJ6qfkmOXy2C; reg [2:0] i2IIQfdSjOGJ0HAlaZdYe; reg [1:0] xSW8arCNXsyV5zIEXuGUQB; reg [1:0] ck9Ya76HU61qWvvl3qwfRG; reg [2:0] dQhJtS5aSGZCPWaJqkkHi; reg t69iUVjqBKXZw2tNuE5YceG; reg [1:0] BNI9VucWF1TWsCAM4sBCHE; reg EIfu64RX7LMQGnynQeCGuD; reg [2:0] KlzCAte3JMaaOEkO4JjiQD; reg adAAE3kEND2Qg9vtBb6GhC; reg RDHFrcFHrfEJ7yzR8LWzB; reg m9VM4i4cuk6jpZ1rsm5lI2C; wire UQZu8I6cZaXNq9rOGDXlJF; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : h6oTzWU1a3otHwaiji95ID if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin JomiEQo6ylRrlhLJPFsQTG <= 3'b000; GP01IUV0xObQQCSdqL463C <= 3'b000; X7FJ0jgk6hqdMN8BingGvE <= 2'b00; WXS42gmgDxS46057b3AGD <= 2'b00; mb13NdjIe7rpJDLNih8AaE <= 2'b00; pDYTWTp6fyrEdA1XnDiP6E <= 1'b0; Xf88wK4mkniJ6qfkmOXy2C <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin JomiEQo6ylRrlhLJPFsQTG <= 3'b000; GP01IUV0xObQQCSdqL463C <= 3'b000; X7FJ0jgk6hqdMN8BingGvE <= 2'b00; WXS42gmgDxS46057b3AGD <= 2'b00; mb13NdjIe7rpJDLNih8AaE <= 2'b00; pDYTWTp6fyrEdA1XnDiP6E <= 1'b0; Xf88wK4mkniJ6qfkmOXy2C <= 1'b0; end else begin JomiEQo6ylRrlhLJPFsQTG <= i2IIQfdSjOGJ0HAlaZdYe; X7FJ0jgk6hqdMN8BingGvE <= xSW8arCNXsyV5zIEXuGUQB; WXS42gmgDxS46057b3AGD <= ck9Ya76HU61qWvvl3qwfRG; GP01IUV0xObQQCSdqL463C <= dQhJtS5aSGZCPWaJqkkHi; pDYTWTp6fyrEdA1XnDiP6E <= t69iUVjqBKXZw2tNuE5YceG; mb13NdjIe7rpJDLNih8AaE <= BNI9VucWF1TWsCAM4sBCHE; Xf88wK4mkniJ6qfkmOXy2C <= EIfu64RX7LMQGnynQeCGuD; end end end always @(Ck459KQ1C8vRbine3lrkt, DCqZJgzh8RI4wgf1TYRoc, GP01IUV0xObQQCSdqL463C, JomiEQo6ylRrlhLJPFsQTG, WXS42gmgDxS46057b3AGD, X7FJ0jgk6hqdMN8BingGvE, Xf88wK4mkniJ6qfkmOXy2C, mb13NdjIe7rpJDLNih8AaE, pDYTWTp6fyrEdA1XnDiP6E) begin i2IIQfdSjOGJ0HAlaZdYe = JomiEQo6ylRrlhLJPFsQTG; xSW8arCNXsyV5zIEXuGUQB = X7FJ0jgk6hqdMN8BingGvE; ck9Ya76HU61qWvvl3qwfRG = WXS42gmgDxS46057b3AGD; dQhJtS5aSGZCPWaJqkkHi = GP01IUV0xObQQCSdqL463C; t69iUVjqBKXZw2tNuE5YceG = pDYTWTp6fyrEdA1XnDiP6E; BNI9VucWF1TWsCAM4sBCHE = mb13NdjIe7rpJDLNih8AaE; EIfu64RX7LMQGnynQeCGuD = Xf88wK4mkniJ6qfkmOXy2C; case ( mb13NdjIe7rpJDLNih8AaE) 2'b00 : begin BNI9VucWF1TWsCAM4sBCHE = 2'b00; EIfu64RX7LMQGnynQeCGuD = 1'b0; if (WXS42gmgDxS46057b3AGD == 2'b01) begin BNI9VucWF1TWsCAM4sBCHE = 2'b01; end end 2'b01 : begin EIfu64RX7LMQGnynQeCGuD = ! (GP01IUV0xObQQCSdqL463C <= 3'b011); if (WXS42gmgDxS46057b3AGD == 2'b10) begin BNI9VucWF1TWsCAM4sBCHE = 2'b10; end end 2'b10 : begin EIfu64RX7LMQGnynQeCGuD = 1'b0; if (WXS42gmgDxS46057b3AGD == 2'b01) begin BNI9VucWF1TWsCAM4sBCHE = 2'b11; end end 2'b11 : begin if (WXS42gmgDxS46057b3AGD == 2'b01) begin BNI9VucWF1TWsCAM4sBCHE = 2'b11; EIfu64RX7LMQGnynQeCGuD = ! (GP01IUV0xObQQCSdqL463C <= 3'b011); end else begin EIfu64RX7LMQGnynQeCGuD = 1'b0; BNI9VucWF1TWsCAM4sBCHE = 2'b00; end end default : begin BNI9VucWF1TWsCAM4sBCHE = 2'b00; EIfu64RX7LMQGnynQeCGuD = 1'b0; end endcase case ( WXS42gmgDxS46057b3AGD) 2'b00 : begin ck9Ya76HU61qWvvl3qwfRG = 2'b00; dQhJtS5aSGZCPWaJqkkHi = 3'b000; adAAE3kEND2Qg9vtBb6GhC = 1'b0; if (Ck459KQ1C8vRbine3lrkt && (JomiEQo6ylRrlhLJPFsQTG == 3'b111)) begin ck9Ya76HU61qWvvl3qwfRG = 2'b01; end end 2'b01 : begin ck9Ya76HU61qWvvl3qwfRG = 2'b01; adAAE3kEND2Qg9vtBb6GhC = DCqZJgzh8RI4wgf1TYRoc; if (DCqZJgzh8RI4wgf1TYRoc) begin if (GP01IUV0xObQQCSdqL463C == 3'b111) begin ck9Ya76HU61qWvvl3qwfRG = 2'b10; end dQhJtS5aSGZCPWaJqkkHi = GP01IUV0xObQQCSdqL463C + 3'b001; end end 2'b10 : begin adAAE3kEND2Qg9vtBb6GhC = 1'b0; if (GP01IUV0xObQQCSdqL463C == 3'b111) begin if (Ck459KQ1C8vRbine3lrkt && (JomiEQo6ylRrlhLJPFsQTG == 3'b111)) begin ck9Ya76HU61qWvvl3qwfRG = 2'b01; end else begin ck9Ya76HU61qWvvl3qwfRG = 2'b00; end end dQhJtS5aSGZCPWaJqkkHi = GP01IUV0xObQQCSdqL463C + 3'b001; end default : begin ck9Ya76HU61qWvvl3qwfRG = 2'b00; dQhJtS5aSGZCPWaJqkkHi = 3'b000; adAAE3kEND2Qg9vtBb6GhC = 1'b0; end endcase case ( X7FJ0jgk6hqdMN8BingGvE) 2'b00 : begin xSW8arCNXsyV5zIEXuGUQB = 2'b00; i2IIQfdSjOGJ0HAlaZdYe = 3'b000; t69iUVjqBKXZw2tNuE5YceG = 1'b0; if (Ck459KQ1C8vRbine3lrkt) begin xSW8arCNXsyV5zIEXuGUQB = 2'b01; i2IIQfdSjOGJ0HAlaZdYe = 3'b001; end end 2'b01 : begin xSW8arCNXsyV5zIEXuGUQB = 2'b01; t69iUVjqBKXZw2tNuE5YceG = 1'b0; if (Ck459KQ1C8vRbine3lrkt) begin if (JomiEQo6ylRrlhLJPFsQTG == 3'b111) begin xSW8arCNXsyV5zIEXuGUQB = 2'b10; t69iUVjqBKXZw2tNuE5YceG = 1'b1; end else begin xSW8arCNXsyV5zIEXuGUQB = 2'b01; end i2IIQfdSjOGJ0HAlaZdYe = JomiEQo6ylRrlhLJPFsQTG + 3'b001; end end 2'b10 : begin xSW8arCNXsyV5zIEXuGUQB = 2'b10; if (Ck459KQ1C8vRbine3lrkt) begin if (JomiEQo6ylRrlhLJPFsQTG == 3'b111) begin xSW8arCNXsyV5zIEXuGUQB = 2'b01; t69iUVjqBKXZw2tNuE5YceG = 1'b0; end else begin xSW8arCNXsyV5zIEXuGUQB = 2'b10; t69iUVjqBKXZw2tNuE5YceG = 1'b1; end i2IIQfdSjOGJ0HAlaZdYe = JomiEQo6ylRrlhLJPFsQTG + 3'b001; end end default : begin xSW8arCNXsyV5zIEXuGUQB = 2'b00; i2IIQfdSjOGJ0HAlaZdYe = 3'b111; t69iUVjqBKXZw2tNuE5YceG = 1'b0; end endcase KlzCAte3JMaaOEkO4JjiQD = GP01IUV0xObQQCSdqL463C; RDHFrcFHrfEJ7yzR8LWzB = pDYTWTp6fyrEdA1XnDiP6E; m9VM4i4cuk6jpZ1rsm5lI2C = Xf88wK4mkniJ6qfkmOXy2C; end assign MCqIdNMOB0Mg1cefHLMjpH = KlzCAte3JMaaOEkO4JjiQD; assign j41GwwL8b9NI9l6ZScQ1PbG = adAAE3kEND2Qg9vtBb6GhC; assign i8H7HzN3cvjFks6MZ5qaqF = RDHFrcFHrfEJ7yzR8LWzB; assign SAcShGLK2YZQrWHGqGVvjD = m9VM4i4cuk6jpZ1rsm5lI2C; endmodule