`timescale 1 ns / 1 ns module HMcgSDBQI8srN5Fet9wEnG (v04pHKxyc2sPW047bbyUgE, JAMOfrNHxGSYDF0urqkLN, NHkD6RGVcC6B7ibmcHypOC, n6CG7K4rgMGw86VJoKnfuOD, R6zf5iqRNVEGVBO8egq8kF, u6oVvmCf0f079jLPodlV5B, qv4pS1KBm1VYTuOTZHo04F, LSv5mOYTPLq5vaIpiVTypC); input v04pHKxyc2sPW047bbyUgE; input JAMOfrNHxGSYDF0urqkLN; input NHkD6RGVcC6B7ibmcHypOC; input n6CG7K4rgMGw86VJoKnfuOD; input R6zf5iqRNVEGVBO8egq8kF; output [1:0] u6oVvmCf0f079jLPodlV5B; output qv4pS1KBm1VYTuOTZHo04F; output LSv5mOYTPLq5vaIpiVTypC; reg [1:0] JomiEQo6ylRrlhLJPFsQTG; reg [1:0] X7FJ0jgk6hqdMN8BingGvE; reg [1:0] WXS42gmgDxS46057b3AGD; reg [1:0] GP01IUV0xObQQCSdqL463C; reg pDYTWTp6fyrEdA1XnDiP6E; reg [1:0] mb13NdjIe7rpJDLNih8AaE; reg Xf88wK4mkniJ6qfkmOXy2C; reg [1:0] i2IIQfdSjOGJ0HAlaZdYe; reg [1:0] xSW8arCNXsyV5zIEXuGUQB; reg [1:0] ck9Ya76HU61qWvvl3qwfRG; reg [1:0] dQhJtS5aSGZCPWaJqkkHi; reg t69iUVjqBKXZw2tNuE5YceG; reg [1:0] BNI9VucWF1TWsCAM4sBCHE; reg EIfu64RX7LMQGnynQeCGuD; reg [1:0] kQTKPzorXSE4AAa1J1hLMC; reg pOtk3FXvlf4GjzqBlLmJ; reg p1eTMzAax3btlf0uh4lGPB; reg vowCHQiasjCt8aFj2iOmDC; wire PPqzwNg6rSKimNIAzt6NoB; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : h6oTzWU1a3otHwaiji95ID if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin JomiEQo6ylRrlhLJPFsQTG <= 2'b00; GP01IUV0xObQQCSdqL463C <= 2'b00; X7FJ0jgk6hqdMN8BingGvE <= 2'b00; WXS42gmgDxS46057b3AGD <= 2'b00; mb13NdjIe7rpJDLNih8AaE <= 2'b00; pDYTWTp6fyrEdA1XnDiP6E <= 1'b0; Xf88wK4mkniJ6qfkmOXy2C <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin JomiEQo6ylRrlhLJPFsQTG <= 2'b00; GP01IUV0xObQQCSdqL463C <= 2'b00; X7FJ0jgk6hqdMN8BingGvE <= 2'b00; WXS42gmgDxS46057b3AGD <= 2'b00; mb13NdjIe7rpJDLNih8AaE <= 2'b00; pDYTWTp6fyrEdA1XnDiP6E <= 1'b0; Xf88wK4mkniJ6qfkmOXy2C <= 1'b0; end else begin JomiEQo6ylRrlhLJPFsQTG <= i2IIQfdSjOGJ0HAlaZdYe; X7FJ0jgk6hqdMN8BingGvE <= xSW8arCNXsyV5zIEXuGUQB; WXS42gmgDxS46057b3AGD <= ck9Ya76HU61qWvvl3qwfRG; GP01IUV0xObQQCSdqL463C <= dQhJtS5aSGZCPWaJqkkHi; pDYTWTp6fyrEdA1XnDiP6E <= t69iUVjqBKXZw2tNuE5YceG; mb13NdjIe7rpJDLNih8AaE <= BNI9VucWF1TWsCAM4sBCHE; Xf88wK4mkniJ6qfkmOXy2C <= EIfu64RX7LMQGnynQeCGuD; end end end always @(GP01IUV0xObQQCSdqL463C, JomiEQo6ylRrlhLJPFsQTG, NHkD6RGVcC6B7ibmcHypOC, WXS42gmgDxS46057b3AGD, X7FJ0jgk6hqdMN8BingGvE, Xf88wK4mkniJ6qfkmOXy2C, mb13NdjIe7rpJDLNih8AaE, n6CG7K4rgMGw86VJoKnfuOD, pDYTWTp6fyrEdA1XnDiP6E) begin i2IIQfdSjOGJ0HAlaZdYe = JomiEQo6ylRrlhLJPFsQTG; xSW8arCNXsyV5zIEXuGUQB = X7FJ0jgk6hqdMN8BingGvE; ck9Ya76HU61qWvvl3qwfRG = WXS42gmgDxS46057b3AGD; dQhJtS5aSGZCPWaJqkkHi = GP01IUV0xObQQCSdqL463C; t69iUVjqBKXZw2tNuE5YceG = pDYTWTp6fyrEdA1XnDiP6E; BNI9VucWF1TWsCAM4sBCHE = mb13NdjIe7rpJDLNih8AaE; EIfu64RX7LMQGnynQeCGuD = Xf88wK4mkniJ6qfkmOXy2C; case ( mb13NdjIe7rpJDLNih8AaE) 2'b00 : begin BNI9VucWF1TWsCAM4sBCHE = 2'b00; EIfu64RX7LMQGnynQeCGuD = 1'b0; if (WXS42gmgDxS46057b3AGD == 2'b01) begin BNI9VucWF1TWsCAM4sBCHE = 2'b01; end end 2'b01 : begin EIfu64RX7LMQGnynQeCGuD = ! (GP01IUV0xObQQCSdqL463C <= 2'b01); if (WXS42gmgDxS46057b3AGD == 2'b10) begin BNI9VucWF1TWsCAM4sBCHE = 2'b10; end end 2'b10 : begin EIfu64RX7LMQGnynQeCGuD = 1'b0; if (WXS42gmgDxS46057b3AGD == 2'b01) begin BNI9VucWF1TWsCAM4sBCHE = 2'b11; end end 2'b11 : begin if (WXS42gmgDxS46057b3AGD == 2'b01) begin BNI9VucWF1TWsCAM4sBCHE = 2'b11; EIfu64RX7LMQGnynQeCGuD = ! (GP01IUV0xObQQCSdqL463C <= 2'b01); end else begin EIfu64RX7LMQGnynQeCGuD = 1'b0; BNI9VucWF1TWsCAM4sBCHE = 2'b00; end end default : begin BNI9VucWF1TWsCAM4sBCHE = 2'b00; EIfu64RX7LMQGnynQeCGuD = 1'b0; end endcase case ( WXS42gmgDxS46057b3AGD) 2'b00 : begin ck9Ya76HU61qWvvl3qwfRG = 2'b00; dQhJtS5aSGZCPWaJqkkHi = 2'b00; pOtk3FXvlf4GjzqBlLmJ = 1'b0; if (NHkD6RGVcC6B7ibmcHypOC && (JomiEQo6ylRrlhLJPFsQTG == 2'b11)) begin ck9Ya76HU61qWvvl3qwfRG = 2'b01; end end 2'b01 : begin ck9Ya76HU61qWvvl3qwfRG = 2'b01; pOtk3FXvlf4GjzqBlLmJ = n6CG7K4rgMGw86VJoKnfuOD; if (n6CG7K4rgMGw86VJoKnfuOD) begin if (GP01IUV0xObQQCSdqL463C == 2'b11) begin ck9Ya76HU61qWvvl3qwfRG = 2'b10; end dQhJtS5aSGZCPWaJqkkHi = GP01IUV0xObQQCSdqL463C + 2'b01; end end 2'b10 : begin pOtk3FXvlf4GjzqBlLmJ = 1'b0; if (GP01IUV0xObQQCSdqL463C == 2'b11) begin if (NHkD6RGVcC6B7ibmcHypOC && (JomiEQo6ylRrlhLJPFsQTG == 2'b11)) begin ck9Ya76HU61qWvvl3qwfRG = 2'b01; end else begin ck9Ya76HU61qWvvl3qwfRG = 2'b00; end end dQhJtS5aSGZCPWaJqkkHi = GP01IUV0xObQQCSdqL463C + 2'b01; end default : begin ck9Ya76HU61qWvvl3qwfRG = 2'b00; dQhJtS5aSGZCPWaJqkkHi = 2'b00; pOtk3FXvlf4GjzqBlLmJ = 1'b0; end endcase case ( X7FJ0jgk6hqdMN8BingGvE) 2'b00 : begin xSW8arCNXsyV5zIEXuGUQB = 2'b00; i2IIQfdSjOGJ0HAlaZdYe = 2'b00; t69iUVjqBKXZw2tNuE5YceG = 1'b0; if (NHkD6RGVcC6B7ibmcHypOC) begin xSW8arCNXsyV5zIEXuGUQB = 2'b01; i2IIQfdSjOGJ0HAlaZdYe = 2'b01; end end 2'b01 : begin xSW8arCNXsyV5zIEXuGUQB = 2'b01; t69iUVjqBKXZw2tNuE5YceG = 1'b0; if (NHkD6RGVcC6B7ibmcHypOC) begin if (JomiEQo6ylRrlhLJPFsQTG == 2'b11) begin xSW8arCNXsyV5zIEXuGUQB = 2'b10; t69iUVjqBKXZw2tNuE5YceG = 1'b1; end else begin xSW8arCNXsyV5zIEXuGUQB = 2'b01; end i2IIQfdSjOGJ0HAlaZdYe = JomiEQo6ylRrlhLJPFsQTG + 2'b01; end end 2'b10 : begin xSW8arCNXsyV5zIEXuGUQB = 2'b10; if (NHkD6RGVcC6B7ibmcHypOC) begin if (JomiEQo6ylRrlhLJPFsQTG == 2'b11) begin xSW8arCNXsyV5zIEXuGUQB = 2'b01; t69iUVjqBKXZw2tNuE5YceG = 1'b0; end else begin xSW8arCNXsyV5zIEXuGUQB = 2'b10; t69iUVjqBKXZw2tNuE5YceG = 1'b1; end i2IIQfdSjOGJ0HAlaZdYe = JomiEQo6ylRrlhLJPFsQTG + 2'b01; end end default : begin xSW8arCNXsyV5zIEXuGUQB = 2'b00; i2IIQfdSjOGJ0HAlaZdYe = 2'b11; t69iUVjqBKXZw2tNuE5YceG = 1'b0; end endcase kQTKPzorXSE4AAa1J1hLMC = GP01IUV0xObQQCSdqL463C; p1eTMzAax3btlf0uh4lGPB = pDYTWTp6fyrEdA1XnDiP6E; vowCHQiasjCt8aFj2iOmDC = Xf88wK4mkniJ6qfkmOXy2C; end assign u6oVvmCf0f079jLPodlV5B = kQTKPzorXSE4AAa1J1hLMC; assign qv4pS1KBm1VYTuOTZHo04F = pOtk3FXvlf4GjzqBlLmJ; assign LSv5mOYTPLq5vaIpiVTypC = p1eTMzAax3btlf0uh4lGPB; endmodule