`timescale 1 ns / 1 ns module QCP2KsVCXOv9pucMwLlsBG (tu9ohhJdK00us7wfvWNQYC, utKZyKAnyhCUOZ6LUagX4D, gA7z08sAKJH0Dq3fae8ZeF, vrNoBb2ZnRj9xKaojUq7EG, IS0z2hJ2LtWljhJ4YYLYaE, TkIATgh1a29iglca8RarC, b4TwkCZxxInAgelXDhMy8E, f9IpN1esn9PJkU40eAffHB, ySOrNaQmYucOX4cyOT5LnG, gmoWrkWFJMiyePfRw5V1lD, nzbLrBOekdX928cLtCU5jD, a9DSedGWFdieeZlu7mhtF7D, zzBKVZ6VX4ht5u9x9EjCiD, j83GXtGY1eMU252JJ6B9mC, r7Q5mFJeRMLiOPMHQDcQQB, wtshVXYU5akP8bsJW8meZH, w2g8aZ7DNLiB7xd9ema9tID, EpypH5ZIz8rvw2qkajrEUD, k5yT5mPpUVKMKN3fkRm1LR, hfxEgMPHtdNs5za4aJfZR); input signed [32:0] tu9ohhJdK00us7wfvWNQYC; input signed [32:0] utKZyKAnyhCUOZ6LUagX4D; input signed [32:0] gA7z08sAKJH0Dq3fae8ZeF; input signed [32:0] vrNoBb2ZnRj9xKaojUq7EG; input signed [15:0] IS0z2hJ2LtWljhJ4YYLYaE; input signed [15:0] TkIATgh1a29iglca8RarC; input signed [15:0] b4TwkCZxxInAgelXDhMy8E; input signed [15:0] f9IpN1esn9PJkU40eAffHB; input signed [15:0] ySOrNaQmYucOX4cyOT5LnG; input signed [15:0] gmoWrkWFJMiyePfRw5V1lD; input signed [15:0] nzbLrBOekdX928cLtCU5jD; input signed [15:0] a9DSedGWFdieeZlu7mhtF7D; output signed [15:0] zzBKVZ6VX4ht5u9x9EjCiD; output signed [15:0] j83GXtGY1eMU252JJ6B9mC; output signed [15:0] r7Q5mFJeRMLiOPMHQDcQQB; output signed [15:0] wtshVXYU5akP8bsJW8meZH; output signed [15:0] w2g8aZ7DNLiB7xd9ema9tID; output signed [15:0] EpypH5ZIz8rvw2qkajrEUD; output signed [15:0] k5yT5mPpUVKMKN3fkRm1LR; output signed [15:0] hfxEgMPHtdNs5za4aJfZR; wire signed [15:0] NepiOXZuBICFGpeGQlYktD [0:3]; wire signed [15:0] UXv2GwCr4OuG2xYfnBhfl [0:3]; wire signed [15:0] T32N7tx3lM4AhPeUl37rcH; wire signed [15:0] gfHKuOgIEm3NEBVOtR9xpG; wire signed [15:0] hHN5I2JoMoPUhhDXhbQxrC; wire signed [15:0] w79PUgPPTaX91btJC6rBPH; wire signed [15:0] HjSWL8FbBbt7xPnQaMIEbF; wire signed [15:0] f7F3bB4hbBp3mLhQVQqnlGC; wire signed [15:0] c0BcY26HQrpNGiwSIvA5UWF; wire signed [15:0] Vrc585EEynXhU8ctzsDNfH; wire BsfHWou9QgD6rZmrYrQfXG; assign NepiOXZuBICFGpeGQlYktD[0] = IS0z2hJ2LtWljhJ4YYLYaE; assign NepiOXZuBICFGpeGQlYktD[1] = TkIATgh1a29iglca8RarC; assign NepiOXZuBICFGpeGQlYktD[2] = b4TwkCZxxInAgelXDhMy8E; assign NepiOXZuBICFGpeGQlYktD[3] = f9IpN1esn9PJkU40eAffHB; assign UXv2GwCr4OuG2xYfnBhfl[0] = ySOrNaQmYucOX4cyOT5LnG; assign UXv2GwCr4OuG2xYfnBhfl[1] = gmoWrkWFJMiyePfRw5V1lD; assign UXv2GwCr4OuG2xYfnBhfl[2] = nzbLrBOekdX928cLtCU5jD; assign UXv2GwCr4OuG2xYfnBhfl[3] = a9DSedGWFdieeZlu7mhtF7D; assign T32N7tx3lM4AhPeUl37rcH = (tu9ohhJdK00us7wfvWNQYC == 33'sh000000000 ? NepiOXZuBICFGpeGQlYktD[0] : (tu9ohhJdK00us7wfvWNQYC == 33'sh000000001 ? NepiOXZuBICFGpeGQlYktD[1] : (tu9ohhJdK00us7wfvWNQYC == 33'sh000000002 ? NepiOXZuBICFGpeGQlYktD[2] : NepiOXZuBICFGpeGQlYktD[3]))); assign gfHKuOgIEm3NEBVOtR9xpG = (tu9ohhJdK00us7wfvWNQYC == 33'sh000000000 ? UXv2GwCr4OuG2xYfnBhfl[0] : (tu9ohhJdK00us7wfvWNQYC == 33'sh000000001 ? UXv2GwCr4OuG2xYfnBhfl[1] : (tu9ohhJdK00us7wfvWNQYC == 33'sh000000002 ? UXv2GwCr4OuG2xYfnBhfl[2] : UXv2GwCr4OuG2xYfnBhfl[3]))); assign zzBKVZ6VX4ht5u9x9EjCiD = T32N7tx3lM4AhPeUl37rcH; assign hHN5I2JoMoPUhhDXhbQxrC = (utKZyKAnyhCUOZ6LUagX4D == 33'sh000000000 ? NepiOXZuBICFGpeGQlYktD[0] : (utKZyKAnyhCUOZ6LUagX4D == 33'sh000000001 ? NepiOXZuBICFGpeGQlYktD[1] : (utKZyKAnyhCUOZ6LUagX4D == 33'sh000000002 ? NepiOXZuBICFGpeGQlYktD[2] : NepiOXZuBICFGpeGQlYktD[3]))); assign w79PUgPPTaX91btJC6rBPH = (utKZyKAnyhCUOZ6LUagX4D == 33'sh000000000 ? UXv2GwCr4OuG2xYfnBhfl[0] : (utKZyKAnyhCUOZ6LUagX4D == 33'sh000000001 ? UXv2GwCr4OuG2xYfnBhfl[1] : (utKZyKAnyhCUOZ6LUagX4D == 33'sh000000002 ? UXv2GwCr4OuG2xYfnBhfl[2] : UXv2GwCr4OuG2xYfnBhfl[3]))); assign j83GXtGY1eMU252JJ6B9mC = hHN5I2JoMoPUhhDXhbQxrC; assign HjSWL8FbBbt7xPnQaMIEbF = (gA7z08sAKJH0Dq3fae8ZeF == 33'sh000000000 ? NepiOXZuBICFGpeGQlYktD[0] : (gA7z08sAKJH0Dq3fae8ZeF == 33'sh000000001 ? NepiOXZuBICFGpeGQlYktD[1] : (gA7z08sAKJH0Dq3fae8ZeF == 33'sh000000002 ? NepiOXZuBICFGpeGQlYktD[2] : NepiOXZuBICFGpeGQlYktD[3]))); assign f7F3bB4hbBp3mLhQVQqnlGC = (gA7z08sAKJH0Dq3fae8ZeF == 33'sh000000000 ? UXv2GwCr4OuG2xYfnBhfl[0] : (gA7z08sAKJH0Dq3fae8ZeF == 33'sh000000001 ? UXv2GwCr4OuG2xYfnBhfl[1] : (gA7z08sAKJH0Dq3fae8ZeF == 33'sh000000002 ? UXv2GwCr4OuG2xYfnBhfl[2] : UXv2GwCr4OuG2xYfnBhfl[3]))); assign r7Q5mFJeRMLiOPMHQDcQQB = HjSWL8FbBbt7xPnQaMIEbF; assign c0BcY26HQrpNGiwSIvA5UWF = (vrNoBb2ZnRj9xKaojUq7EG == 33'sh000000000 ? NepiOXZuBICFGpeGQlYktD[0] : (vrNoBb2ZnRj9xKaojUq7EG == 33'sh000000001 ? NepiOXZuBICFGpeGQlYktD[1] : (vrNoBb2ZnRj9xKaojUq7EG == 33'sh000000002 ? NepiOXZuBICFGpeGQlYktD[2] : NepiOXZuBICFGpeGQlYktD[3]))); assign Vrc585EEynXhU8ctzsDNfH = (vrNoBb2ZnRj9xKaojUq7EG == 33'sh000000000 ? UXv2GwCr4OuG2xYfnBhfl[0] : (vrNoBb2ZnRj9xKaojUq7EG == 33'sh000000001 ? UXv2GwCr4OuG2xYfnBhfl[1] : (vrNoBb2ZnRj9xKaojUq7EG == 33'sh000000002 ? UXv2GwCr4OuG2xYfnBhfl[2] : UXv2GwCr4OuG2xYfnBhfl[3]))); assign wtshVXYU5akP8bsJW8meZH = c0BcY26HQrpNGiwSIvA5UWF; assign w2g8aZ7DNLiB7xd9ema9tID = gfHKuOgIEm3NEBVOtR9xpG; assign EpypH5ZIz8rvw2qkajrEUD = w79PUgPPTaX91btJC6rBPH; assign k5yT5mPpUVKMKN3fkRm1LR = f7F3bB4hbBp3mLhQVQqnlGC; assign hfxEgMPHtdNs5za4aJfZR = Vrc585EEynXhU8ctzsDNfH; endmodule