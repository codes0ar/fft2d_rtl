`timescale 1 ns / 1 ns module CF4YZpD8T3bZDeoOS74nFB (v04pHKxyc2sPW047bbyUgE, JAMOfrNHxGSYDF0urqkLN, kIsHJAwQMWbIiCsXfX1rTG, DKGIysOp4cb2Wy4ifYHB8D, R6zf5iqRNVEGVBO8egq8kF, yTf5WZbZOLm2uKwJmXk5sG, wGlnEfCkRPxniOjCaZH6XG, RDvlVEJspE7WkJvNmR8a6C); input v04pHKxyc2sPW047bbyUgE; input JAMOfrNHxGSYDF0urqkLN; input kIsHJAwQMWbIiCsXfX1rTG; input DKGIysOp4cb2Wy4ifYHB8D; input R6zf5iqRNVEGVBO8egq8kF; output [4:0] yTf5WZbZOLm2uKwJmXk5sG; output wGlnEfCkRPxniOjCaZH6XG; output RDvlVEJspE7WkJvNmR8a6C; reg [4:0] JomiEQo6ylRrlhLJPFsQTG; reg [1:0] X7FJ0jgk6hqdMN8BingGvE; reg [1:0] WXS42gmgDxS46057b3AGD; reg [4:0] GP01IUV0xObQQCSdqL463C; reg pDYTWTp6fyrEdA1XnDiP6E; reg [1:0] mb13NdjIe7rpJDLNih8AaE; reg Xf88wK4mkniJ6qfkmOXy2C; reg [4:0] i2IIQfdSjOGJ0HAlaZdYe; reg [1:0] xSW8arCNXsyV5zIEXuGUQB; reg [1:0] ck9Ya76HU61qWvvl3qwfRG; reg [4:0] dQhJtS5aSGZCPWaJqkkHi; reg t69iUVjqBKXZw2tNuE5YceG; reg [1:0] BNI9VucWF1TWsCAM4sBCHE; reg EIfu64RX7LMQGnynQeCGuD; reg [4:0] f0LoJaVTftOyaXbKcYjRST; reg udLm1gCfK1bsBCzyYOebLD; reg mjQQDV7qVUmtyjMgSHu2bC; reg S86yDRz3lzvCeFmkKizFJD; wire mIpum4UZCGRlyCDXdGl1tC; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : h6oTzWU1a3otHwaiji95ID if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin JomiEQo6ylRrlhLJPFsQTG <= 5'b00000; GP01IUV0xObQQCSdqL463C <= 5'b00000; X7FJ0jgk6hqdMN8BingGvE <= 2'b00; WXS42gmgDxS46057b3AGD <= 2'b00; mb13NdjIe7rpJDLNih8AaE <= 2'b00; pDYTWTp6fyrEdA1XnDiP6E <= 1'b0; Xf88wK4mkniJ6qfkmOXy2C <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin JomiEQo6ylRrlhLJPFsQTG <= 5'b00000; GP01IUV0xObQQCSdqL463C <= 5'b00000; X7FJ0jgk6hqdMN8BingGvE <= 2'b00; WXS42gmgDxS46057b3AGD <= 2'b00; mb13NdjIe7rpJDLNih8AaE <= 2'b00; pDYTWTp6fyrEdA1XnDiP6E <= 1'b0; Xf88wK4mkniJ6qfkmOXy2C <= 1'b0; end else begin JomiEQo6ylRrlhLJPFsQTG <= i2IIQfdSjOGJ0HAlaZdYe; X7FJ0jgk6hqdMN8BingGvE <= xSW8arCNXsyV5zIEXuGUQB; WXS42gmgDxS46057b3AGD <= ck9Ya76HU61qWvvl3qwfRG; GP01IUV0xObQQCSdqL463C <= dQhJtS5aSGZCPWaJqkkHi; pDYTWTp6fyrEdA1XnDiP6E <= t69iUVjqBKXZw2tNuE5YceG; mb13NdjIe7rpJDLNih8AaE <= BNI9VucWF1TWsCAM4sBCHE; Xf88wK4mkniJ6qfkmOXy2C <= EIfu64RX7LMQGnynQeCGuD; end end end always @(DKGIysOp4cb2Wy4ifYHB8D, GP01IUV0xObQQCSdqL463C, JomiEQo6ylRrlhLJPFsQTG, WXS42gmgDxS46057b3AGD, X7FJ0jgk6hqdMN8BingGvE, Xf88wK4mkniJ6qfkmOXy2C, kIsHJAwQMWbIiCsXfX1rTG, mb13NdjIe7rpJDLNih8AaE, pDYTWTp6fyrEdA1XnDiP6E) begin i2IIQfdSjOGJ0HAlaZdYe = JomiEQo6ylRrlhLJPFsQTG; xSW8arCNXsyV5zIEXuGUQB = X7FJ0jgk6hqdMN8BingGvE; ck9Ya76HU61qWvvl3qwfRG = WXS42gmgDxS46057b3AGD; dQhJtS5aSGZCPWaJqkkHi = GP01IUV0xObQQCSdqL463C; t69iUVjqBKXZw2tNuE5YceG = pDYTWTp6fyrEdA1XnDiP6E; BNI9VucWF1TWsCAM4sBCHE = mb13NdjIe7rpJDLNih8AaE; EIfu64RX7LMQGnynQeCGuD = Xf88wK4mkniJ6qfkmOXy2C; case ( mb13NdjIe7rpJDLNih8AaE) 2'b00 : begin BNI9VucWF1TWsCAM4sBCHE = 2'b00; EIfu64RX7LMQGnynQeCGuD = 1'b0; if (WXS42gmgDxS46057b3AGD == 2'b01) begin BNI9VucWF1TWsCAM4sBCHE = 2'b01; end end 2'b01 : begin EIfu64RX7LMQGnynQeCGuD = 1'b0; if (WXS42gmgDxS46057b3AGD == 2'b10) begin BNI9VucWF1TWsCAM4sBCHE = 2'b10; end end 2'b10 : begin EIfu64RX7LMQGnynQeCGuD = 1'b0; if (WXS42gmgDxS46057b3AGD == 2'b01) begin BNI9VucWF1TWsCAM4sBCHE = 2'b11; EIfu64RX7LMQGnynQeCGuD = 1'b1; end end 2'b11 : begin if (WXS42gmgDxS46057b3AGD == 2'b01) begin BNI9VucWF1TWsCAM4sBCHE = 2'b11; EIfu64RX7LMQGnynQeCGuD = 1'b1; end else begin EIfu64RX7LMQGnynQeCGuD = 1'b0; BNI9VucWF1TWsCAM4sBCHE = 2'b00; end end default : begin BNI9VucWF1TWsCAM4sBCHE = 2'b00; EIfu64RX7LMQGnynQeCGuD = 1'b0; end endcase case ( WXS42gmgDxS46057b3AGD) 2'b00 : begin ck9Ya76HU61qWvvl3qwfRG = 2'b00; dQhJtS5aSGZCPWaJqkkHi = 5'b00000; udLm1gCfK1bsBCzyYOebLD = 1'b0; if (kIsHJAwQMWbIiCsXfX1rTG && (JomiEQo6ylRrlhLJPFsQTG == 5'b11111)) begin ck9Ya76HU61qWvvl3qwfRG = 2'b01; end end 2'b01 : begin ck9Ya76HU61qWvvl3qwfRG = 2'b01; udLm1gCfK1bsBCzyYOebLD = DKGIysOp4cb2Wy4ifYHB8D; if (DKGIysOp4cb2Wy4ifYHB8D) begin if (GP01IUV0xObQQCSdqL463C == 5'b11111) begin ck9Ya76HU61qWvvl3qwfRG = 2'b10; end dQhJtS5aSGZCPWaJqkkHi = GP01IUV0xObQQCSdqL463C + 5'b00001; end end 2'b10 : begin udLm1gCfK1bsBCzyYOebLD = 1'b1; if (GP01IUV0xObQQCSdqL463C == 5'b11111) begin if (kIsHJAwQMWbIiCsXfX1rTG && (JomiEQo6ylRrlhLJPFsQTG == 5'b11111)) begin ck9Ya76HU61qWvvl3qwfRG = 2'b01; end else begin ck9Ya76HU61qWvvl3qwfRG = 2'b00; end end dQhJtS5aSGZCPWaJqkkHi = GP01IUV0xObQQCSdqL463C + 5'b00001; end default : begin ck9Ya76HU61qWvvl3qwfRG = 2'b00; dQhJtS5aSGZCPWaJqkkHi = 5'b00000; udLm1gCfK1bsBCzyYOebLD = 1'b0; end endcase case ( X7FJ0jgk6hqdMN8BingGvE) 2'b00 : begin xSW8arCNXsyV5zIEXuGUQB = 2'b00; i2IIQfdSjOGJ0HAlaZdYe = 5'b00000; t69iUVjqBKXZw2tNuE5YceG = 1'b0; if (kIsHJAwQMWbIiCsXfX1rTG) begin xSW8arCNXsyV5zIEXuGUQB = 2'b01; i2IIQfdSjOGJ0HAlaZdYe = 5'b00001; end end 2'b01 : begin xSW8arCNXsyV5zIEXuGUQB = 2'b01; t69iUVjqBKXZw2tNuE5YceG = 1'b0; if (kIsHJAwQMWbIiCsXfX1rTG) begin if (JomiEQo6ylRrlhLJPFsQTG == 5'b11111) begin xSW8arCNXsyV5zIEXuGUQB = 2'b10; t69iUVjqBKXZw2tNuE5YceG = 1'b1; end else begin xSW8arCNXsyV5zIEXuGUQB = 2'b01; end i2IIQfdSjOGJ0HAlaZdYe = JomiEQo6ylRrlhLJPFsQTG + 5'b00001; end end 2'b10 : begin xSW8arCNXsyV5zIEXuGUQB = 2'b10; if (kIsHJAwQMWbIiCsXfX1rTG) begin if (JomiEQo6ylRrlhLJPFsQTG == 5'b11111) begin xSW8arCNXsyV5zIEXuGUQB = 2'b01; t69iUVjqBKXZw2tNuE5YceG = 1'b0; end else begin xSW8arCNXsyV5zIEXuGUQB = 2'b10; t69iUVjqBKXZw2tNuE5YceG = 1'b1; end i2IIQfdSjOGJ0HAlaZdYe = JomiEQo6ylRrlhLJPFsQTG + 5'b00001; end end default : begin xSW8arCNXsyV5zIEXuGUQB = 2'b00; i2IIQfdSjOGJ0HAlaZdYe = 5'b11111; t69iUVjqBKXZw2tNuE5YceG = 1'b0; end endcase f0LoJaVTftOyaXbKcYjRST = GP01IUV0xObQQCSdqL463C; mjQQDV7qVUmtyjMgSHu2bC = pDYTWTp6fyrEdA1XnDiP6E; S86yDRz3lzvCeFmkKizFJD = Xf88wK4mkniJ6qfkmOXy2C; end assign yTf5WZbZOLm2uKwJmXk5sG = f0LoJaVTftOyaXbKcYjRST; assign wGlnEfCkRPxniOjCaZH6XG = udLm1gCfK1bsBCzyYOebLD; assign RDvlVEJspE7WkJvNmR8a6C = mjQQDV7qVUmtyjMgSHu2bC; endmodule