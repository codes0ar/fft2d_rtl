`timescale 1 ns / 1 ns module l9MJ6AwAxJzPDBhrXOVFEiF (v04pHKxyc2sPW047bbyUgE, JAMOfrNHxGSYDF0urqkLN, BXAaMHpKzPpYZGFRqoevNE, czP63K90EaJdtsY9EHZ30D, v6PtMRDEb2KzMpzXWCSiwkB, u6oVvmCf0f079jLPodlV5B, qv4pS1KBm1VYTuOTZHo04F, mxtJaiWQH83FcZ66WqnMiH, MtlWbaE0z2xTCIy368PlWF, LSv5mOYTPLq5vaIpiVTypC, R6zf5iqRNVEGVBO8egq8kF, Sek0doTmbyRuabtHW5JKgH, h4q2yYljVPy2UhMxEpHXfqG); input v04pHKxyc2sPW047bbyUgE; input JAMOfrNHxGSYDF0urqkLN; input signed [15:0] BXAaMHpKzPpYZGFRqoevNE; input signed [15:0] czP63K90EaJdtsY9EHZ30D; input v6PtMRDEb2KzMpzXWCSiwkB; input [1:0] u6oVvmCf0f079jLPodlV5B; input qv4pS1KBm1VYTuOTZHo04F; input signed [15:0] mxtJaiWQH83FcZ66WqnMiH; input signed [15:0] MtlWbaE0z2xTCIy368PlWF; input LSv5mOYTPLq5vaIpiVTypC; input R6zf5iqRNVEGVBO8egq8kF; output signed [15:0] Sek0doTmbyRuabtHW5JKgH; output signed [15:0] h4q2yYljVPy2UhMxEpHXfqG; wire signed [15:0] x3T5ivGGBQbBK8kZOoMj3; wire signed [15:0] cMIOWiDVVCoNgM2IifcBEE; wire V1Qnuj0qcpPu0XC8W9in0D; reg de21duRLbf27relCAO1YZB; wire signed [15:0] iOhy3XYM3su7ndksftfCZG; wire [1:0] AECH0r3KnKo0RJFepDhYUD; wire twcuYIJzeZMBjyHmZ1FZDD; wire signed [15:0] dTkGd8OUQ83dmglc4Bt8vF; wire signed [15:0] N2ZdE4zLlq5uRV4rcE2wdE; wire signed [15:0] csMK1iTp18g0vZYjmk9JZD; reg signed [16:0] wFsaSfYltg6TlrWqY1FyGE; reg signed [16:0] T5BRwctOUS2khp8Rzx4l9; reg signed [16:0] t1ZySna7c411biAKwiSaOlF; reg signed [16:0] d8074IV5GByVrE9OuVeZYRF; reg signed [15:0] P6obz6bve3VygHefrMlpoH; reg signed [15:0] v6DJX4vQF6pzvb2z1TWW9LH; reg RwKtM3ApThsv88D4VvltlD; reg signed [15:0] f6eYgeW0rCfd0LIvc2SGHB; reg signed [15:0] m5VNx3xnw67GgdN5661tXkG; reg signed [15:0] IMsvh2kSL36ZxgH6ovKFz; reg signed [15:0] ZvsdK7IB0VkAxGNAOwtzgD; reg q6XydGshj15r9Fju4CQ2iT; reg KuSB40UBeOqvdWcrRv76OB; wire signed [16:0] kHkm1dHei7pqznzynbBKwE; wire signed [16:0] Oym0ZQxbxCKFQ5X3kAuPi; wire signed [16:0] YIMNIvC4K9LQaGT0TCHkcE; wire signed [16:0] IQG3jvRoS6AY8QAkGyV9b; wire signed [16:0] g4G8R7TlPZ9NvGqBSUmdb7F; wire signed [16:0] ndTxZ4yEyGpSsXjLwP10HB; wire signed [16:0] plZaC1IiHJbFqqHndxJpKC; wire signed [16:0] B8fYUIF4y2YvoVPCpuCb0; wire signed [16:0] Yb4qpWQhiQpsJ5laLdw1dG; wire signed [16:0] XETUnhSmrTZNec4mfH5bhE; wire signed [16:0] krcDen5cyZ3crTZ2yfXap; wire signed [16:0] fpzEAgYwqhsLsJYv4qlk8E; wire signed [16:0] n0J4kP9YDHfDkhTNLn56dJ; wire signed [16:0] UpDw6anZs0bMPETxgXld9F; wire signed [16:0] b31KhkrKeVwOtEcPIkvs3; wire signed [16:0] Lcbc8UkQ7CVMIZTyIGqp7G; wire signed [16:0] KinlMSwCRgZdG2BmpRDJAG; wire signed [16:0] t1uTFhJAosQhy0vBWGPplXD; wire signed [16:0] Pr2dhfiX07pLlRUhRGiSR; wire signed [16:0] LgvxMrXuJRlmlCyhLVJYyE; wire signed [16:0] ATjS2KECQ0ZiH7CL8LEnE; wire signed [16:0] RPKurxOe2f65XPpdjKRZMF; wire signed [16:0] a2Lel9XzXgLNrkI13pSAHKE; wire signed [16:0] VJAT39ZYYYO4RWA7Qqf56F; reg signed [15:0] mgknRxAcgFrHqTt5CZvnSF; reg signed [15:0] sCFM4WicR6deeSAdSwumP; reg BKNY6GzA6oGZumjzTATycD; wire signed [15:0] uUcj3UAzjmPW47yNyzbT8C; wire signed [15:0] uwZv0qzQLi0MDBWLWzKuAG; wire n65LdbEr6NMNaEFcjX8Fh6F; wire signed [15:0] x9j7a5gok64zzNKnvdJNnE; wire signed [15:0] bPL0FcLvoxhO0amTUOV9QC; wire signed [15:0] r4JngA0ZVhEElGRZci9fohF; wire signed [15:0] a8xx20Fc5nKc8DbqSwNBuB; reg vLT6ef7BJliTDpt4k5jqF; wire WV3pqDZm8AvqqMyzDNeP3C; xpufpjE4HLrRCiDyZwJhUH ftPsaxEa6Qv5RNEVVRTJoH (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .BXAaMHpKzPpYZGFRqoevNE(BXAaMHpKzPpYZGFRqoevNE), .czP63K90EaJdtsY9EHZ30D(czP63K90EaJdtsY9EHZ30D), .v6PtMRDEb2KzMpzXWCSiwkB(v6PtMRDEb2KzMpzXWCSiwkB), .mxtJaiWQH83FcZ66WqnMiH(mxtJaiWQH83FcZ66WqnMiH), .MtlWbaE0z2xTCIy368PlWF(MtlWbaE0z2xTCIy368PlWF), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .x3T5ivGGBQbBK8kZOoMj3(x3T5ivGGBQbBK8kZOoMj3), .cMIOWiDVVCoNgM2IifcBEE(cMIOWiDVVCoNgM2IifcBEE), .V1Qnuj0qcpPu0XC8W9in0D(V1Qnuj0qcpPu0XC8W9in0D) ); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : MczQYJ6MT1pYZD7C1UhQv if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin de21duRLbf27relCAO1YZB <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin de21duRLbf27relCAO1YZB <= 1'b0; end else begin de21duRLbf27relCAO1YZB <= qv4pS1KBm1VYTuOTZHo04F; end end end PxGtD8RdpEuqNR1OqCny8D #(.AddrWidth(2), .DataWidth(16) ) AnilHth3KIMkOmTekImDLG (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .E7QNJoK4KvAThVFhUlvl2G(iOhy3XYM3su7ndksftfCZG), .l30d1QakAt61ivcMw8sJQE(AECH0r3KnKo0RJFepDhYUD), .UKo8akspo4h0jsZ6g712NB(twcuYIJzeZMBjyHmZ1FZDD), .EYQG62ys4E6V8lISAdlW1C(u6oVvmCf0f079jLPodlV5B), .HmVcl5yQin7hEovf3bwNG(dTkGd8OUQ83dmglc4Bt8vF) ); PxGtD8RdpEuqNR1OqCny8D #(.AddrWidth(2), .DataWidth(16) ) lP1PwnrYvoFkexN79O1XXH (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .E7QNJoK4KvAThVFhUlvl2G(N2ZdE4zLlq5uRV4rcE2wdE), .l30d1QakAt61ivcMw8sJQE(AECH0r3KnKo0RJFepDhYUD), .UKo8akspo4h0jsZ6g712NB(twcuYIJzeZMBjyHmZ1FZDD), .EYQG62ys4E6V8lISAdlW1C(u6oVvmCf0f079jLPodlV5B), .HmVcl5yQin7hEovf3bwNG(csMK1iTp18g0vZYjmk9JZD) ); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : plVzUyM9ssc0g5eFRKR67 if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin wFsaSfYltg6TlrWqY1FyGE <= 17'sb00000000000000000; T5BRwctOUS2khp8Rzx4l9 <= 17'sb00000000000000000; t1ZySna7c411biAKwiSaOlF <= 17'sb00000000000000000; d8074IV5GByVrE9OuVeZYRF <= 17'sb00000000000000000; P6obz6bve3VygHefrMlpoH <= 16'sb0000000000000000; v6DJX4vQF6pzvb2z1TWW9LH <= 16'sb0000000000000000; RwKtM3ApThsv88D4VvltlD <= 1'b0; mgknRxAcgFrHqTt5CZvnSF <= 16'sb0000000000000000; sCFM4WicR6deeSAdSwumP <= 16'sb0000000000000000; BKNY6GzA6oGZumjzTATycD <= 1'b0; f6eYgeW0rCfd0LIvc2SGHB <= 16'sb0000000000000000; m5VNx3xnw67GgdN5661tXkG <= 16'sb0000000000000000; IMsvh2kSL36ZxgH6ovKFz <= 16'sb0000000000000000; ZvsdK7IB0VkAxGNAOwtzgD <= 16'sb0000000000000000; q6XydGshj15r9Fju4CQ2iT <= 1'b0; KuSB40UBeOqvdWcrRv76OB <= 1'b0; vLT6ef7BJliTDpt4k5jqF <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin wFsaSfYltg6TlrWqY1FyGE <= 17'sb00000000000000000; T5BRwctOUS2khp8Rzx4l9 <= 17'sb00000000000000000; t1ZySna7c411biAKwiSaOlF <= 17'sb00000000000000000; d8074IV5GByVrE9OuVeZYRF <= 17'sb00000000000000000; P6obz6bve3VygHefrMlpoH <= 16'sb0000000000000000; v6DJX4vQF6pzvb2z1TWW9LH <= 16'sb0000000000000000; RwKtM3ApThsv88D4VvltlD <= 1'b0; mgknRxAcgFrHqTt5CZvnSF <= 16'sb0000000000000000; sCFM4WicR6deeSAdSwumP <= 16'sb0000000000000000; BKNY6GzA6oGZumjzTATycD <= 1'b0; f6eYgeW0rCfd0LIvc2SGHB <= 16'sb0000000000000000; m5VNx3xnw67GgdN5661tXkG <= 16'sb0000000000000000; IMsvh2kSL36ZxgH6ovKFz <= 16'sb0000000000000000; ZvsdK7IB0VkAxGNAOwtzgD <= 16'sb0000000000000000; q6XydGshj15r9Fju4CQ2iT <= 1'b0; KuSB40UBeOqvdWcrRv76OB <= 1'b0; vLT6ef7BJliTDpt4k5jqF <= 1'b0; end else begin wFsaSfYltg6TlrWqY1FyGE <= kHkm1dHei7pqznzynbBKwE; T5BRwctOUS2khp8Rzx4l9 <= Oym0ZQxbxCKFQ5X3kAuPi; t1ZySna7c411biAKwiSaOlF <= YIMNIvC4K9LQaGT0TCHkcE; d8074IV5GByVrE9OuVeZYRF <= IQG3jvRoS6AY8QAkGyV9b; mgknRxAcgFrHqTt5CZvnSF <= P6obz6bve3VygHefrMlpoH; sCFM4WicR6deeSAdSwumP <= v6DJX4vQF6pzvb2z1TWW9LH; BKNY6GzA6oGZumjzTATycD <= RwKtM3ApThsv88D4VvltlD; vLT6ef7BJliTDpt4k5jqF <= KuSB40UBeOqvdWcrRv76OB; KuSB40UBeOqvdWcrRv76OB <= q6XydGshj15r9Fju4CQ2iT; IMsvh2kSL36ZxgH6ovKFz <= f6eYgeW0rCfd0LIvc2SGHB; ZvsdK7IB0VkAxGNAOwtzgD <= m5VNx3xnw67GgdN5661tXkG; f6eYgeW0rCfd0LIvc2SGHB <= x3T5ivGGBQbBK8kZOoMj3; m5VNx3xnw67GgdN5661tXkG <= cMIOWiDVVCoNgM2IifcBEE; P6obz6bve3VygHefrMlpoH <= csMK1iTp18g0vZYjmk9JZD; v6DJX4vQF6pzvb2z1TWW9LH <= dTkGd8OUQ83dmglc4Bt8vF; RwKtM3ApThsv88D4VvltlD <= de21duRLbf27relCAO1YZB; q6XydGshj15r9Fju4CQ2iT <= LSv5mOYTPLq5vaIpiVTypC && V1Qnuj0qcpPu0XC8W9in0D; end end end assign n65LdbEr6NMNaEFcjX8Fh6F = ( ! LSv5mOYTPLq5vaIpiVTypC) && V1Qnuj0qcpPu0XC8W9in0D; assign KinlMSwCRgZdG2BmpRDJAG = {P6obz6bve3VygHefrMlpoH[15], P6obz6bve3VygHefrMlpoH}; assign t1uTFhJAosQhy0vBWGPplXD = {IMsvh2kSL36ZxgH6ovKFz[15], IMsvh2kSL36ZxgH6ovKFz}; assign kHkm1dHei7pqznzynbBKwE = KinlMSwCRgZdG2BmpRDJAG + t1uTFhJAosQhy0vBWGPplXD; assign Pr2dhfiX07pLlRUhRGiSR = {P6obz6bve3VygHefrMlpoH[15], P6obz6bve3VygHefrMlpoH}; assign LgvxMrXuJRlmlCyhLVJYyE = {IMsvh2kSL36ZxgH6ovKFz[15], IMsvh2kSL36ZxgH6ovKFz}; assign YIMNIvC4K9LQaGT0TCHkcE = Pr2dhfiX07pLlRUhRGiSR - LgvxMrXuJRlmlCyhLVJYyE; assign ATjS2KECQ0ZiH7CL8LEnE = {v6DJX4vQF6pzvb2z1TWW9LH[15], v6DJX4vQF6pzvb2z1TWW9LH}; assign RPKurxOe2f65XPpdjKRZMF = {ZvsdK7IB0VkAxGNAOwtzgD[15], ZvsdK7IB0VkAxGNAOwtzgD}; assign Oym0ZQxbxCKFQ5X3kAuPi = ATjS2KECQ0ZiH7CL8LEnE + RPKurxOe2f65XPpdjKRZMF; assign a2Lel9XzXgLNrkI13pSAHKE = {v6DJX4vQF6pzvb2z1TWW9LH[15], v6DJX4vQF6pzvb2z1TWW9LH}; assign VJAT39ZYYYO4RWA7Qqf56F = {ZvsdK7IB0VkAxGNAOwtzgD[15], ZvsdK7IB0VkAxGNAOwtzgD}; assign IQG3jvRoS6AY8QAkGyV9b = a2Lel9XzXgLNrkI13pSAHKE - VJAT39ZYYYO4RWA7Qqf56F; assign uUcj3UAzjmPW47yNyzbT8C = x3T5ivGGBQbBK8kZOoMj3; assign uwZv0qzQLi0MDBWLWzKuAG = cMIOWiDVVCoNgM2IifcBEE; assign g4G8R7TlPZ9NvGqBSUmdb7F = ({wFsaSfYltg6TlrWqY1FyGE[16], wFsaSfYltg6TlrWqY1FyGE[16:1]}) + $signed({1'b0, wFsaSfYltg6TlrWqY1FyGE[0]}); assign ndTxZ4yEyGpSsXjLwP10HB = g4G8R7TlPZ9NvGqBSUmdb7F >>> 8'd1; assign plZaC1IiHJbFqqHndxJpKC = {ndTxZ4yEyGpSsXjLwP10HB[15:0], 1'b0}; assign x9j7a5gok64zzNKnvdJNnE = plZaC1IiHJbFqqHndxJpKC[15:0]; assign B8fYUIF4y2YvoVPCpuCb0 = ({T5BRwctOUS2khp8Rzx4l9[16], T5BRwctOUS2khp8Rzx4l9[16:1]}) + $signed({1'b0, T5BRwctOUS2khp8Rzx4l9[0]}); assign Yb4qpWQhiQpsJ5laLdw1dG = B8fYUIF4y2YvoVPCpuCb0 >>> 8'd1; assign XETUnhSmrTZNec4mfH5bhE = {Yb4qpWQhiQpsJ5laLdw1dG[15:0], 1'b0}; assign bPL0FcLvoxhO0amTUOV9QC = XETUnhSmrTZNec4mfH5bhE[15:0]; assign krcDen5cyZ3crTZ2yfXap = ({t1ZySna7c411biAKwiSaOlF[16], t1ZySna7c411biAKwiSaOlF[16:1]}) + $signed({1'b0, t1ZySna7c411biAKwiSaOlF[0]}); assign fpzEAgYwqhsLsJYv4qlk8E = krcDen5cyZ3crTZ2yfXap >>> 8'd1; assign n0J4kP9YDHfDkhTNLn56dJ = {fpzEAgYwqhsLsJYv4qlk8E[15:0], 1'b0}; assign r4JngA0ZVhEElGRZci9fohF = n0J4kP9YDHfDkhTNLn56dJ[15:0]; assign UpDw6anZs0bMPETxgXld9F = ({d8074IV5GByVrE9OuVeZYRF[16], d8074IV5GByVrE9OuVeZYRF[16:1]}) + $signed({1'b0, d8074IV5GByVrE9OuVeZYRF[0]}); assign b31KhkrKeVwOtEcPIkvs3 = UpDw6anZs0bMPETxgXld9F >>> 8'd1; assign Lcbc8UkQ7CVMIZTyIGqp7G = {b31KhkrKeVwOtEcPIkvs3[15:0], 1'b0}; assign a8xx20Fc5nKc8DbqSwNBuB = Lcbc8UkQ7CVMIZTyIGqp7G[15:0]; EWb20Zh4qFGY7CXWFWIrfF RXE5sNatFSMdPgXShrZQ1F (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .v6PtMRDEb2KzMpzXWCSiwkB(v6PtMRDEb2KzMpzXWCSiwkB), .mgknRxAcgFrHqTt5CZvnSF(mgknRxAcgFrHqTt5CZvnSF), .sCFM4WicR6deeSAdSwumP(sCFM4WicR6deeSAdSwumP), .BKNY6GzA6oGZumjzTATycD(BKNY6GzA6oGZumjzTATycD), .uUcj3UAzjmPW47yNyzbT8C(uUcj3UAzjmPW47yNyzbT8C), .uwZv0qzQLi0MDBWLWzKuAG(uwZv0qzQLi0MDBWLWzKuAG), .n65LdbEr6NMNaEFcjX8Fh6F(n65LdbEr6NMNaEFcjX8Fh6F), .x9j7a5gok64zzNKnvdJNnE(x9j7a5gok64zzNKnvdJNnE), .bPL0FcLvoxhO0amTUOV9QC(bPL0FcLvoxhO0amTUOV9QC), .r4JngA0ZVhEElGRZci9fohF(r4JngA0ZVhEElGRZci9fohF), .a8xx20Fc5nKc8DbqSwNBuB(a8xx20Fc5nKc8DbqSwNBuB), .vLT6ef7BJliTDpt4k5jqF(vLT6ef7BJliTDpt4k5jqF), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .N2ZdE4zLlq5uRV4rcE2wdE(N2ZdE4zLlq5uRV4rcE2wdE), .iOhy3XYM3su7ndksftfCZG(iOhy3XYM3su7ndksftfCZG), .AECH0r3KnKo0RJFepDhYUD(AECH0r3KnKo0RJFepDhYUD), .twcuYIJzeZMBjyHmZ1FZDD(twcuYIJzeZMBjyHmZ1FZDD), .Sek0doTmbyRuabtHW5JKgH(Sek0doTmbyRuabtHW5JKgH), .h4q2yYljVPy2UhMxEpHXfqG(h4q2yYljVPy2UhMxEpHXfqG) ); endmodule