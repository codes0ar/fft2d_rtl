`timescale 1 ns / 1 ns module YWcbaK4GTT05DhR2SHpPIG (v04pHKxyc2sPW047bbyUgE, JAMOfrNHxGSYDF0urqkLN, NMWfejbHi1tIjFkylFWDkC, R6zf5iqRNVEGVBO8egq8kF, HXT3YNFExOHI94Xq9VVUBG, EI1r2DTkmcgS5siR9DUFpG); input v04pHKxyc2sPW047bbyUgE; input JAMOfrNHxGSYDF0urqkLN; input NMWfejbHi1tIjFkylFWDkC; input R6zf5iqRNVEGVBO8egq8kF; output signed [15:0] HXT3YNFExOHI94Xq9VVUBG; output signed [15:0] EI1r2DTkmcgS5siR9DUFpG; reg [7:0] TE2s9kaW4jbT2yuidpcUIF; reg [1:0] j9GInQQXHbUGPAy0R0X4BQD; reg [2:0] URO3uEJ9VVi4n2rv5pG4XF; reg [9:0] mevVutOyAH9CPJEBvvvxsF; reg [6:0] Mndh5cWFT2MK7irxEkUgvB; reg DSwbuqNl6si2qBBlHlS4m; reg ADYssd29ifP9Cnqtxk4KFH; reg zUwvjmWVganUujWHX9Ik8G; reg [7:0] vyYw1SbJbcSwGlwsC50cRF; reg [1:0] tHBJR87iWmyApKoUBwoC; reg [2:0] ZXzEhgRyMkDiwOKQ1ZyHtH; reg [9:0] vndcJtBZasetzBa7iOZamH; reg [6:0] W3LV4fQGt3vLDwUnzRRUwH; reg t96JNxh4AbzBXPo2zT29dlG; reg ARo3kgZ8gBa9Exsckya1UB; reg IvvfGB2My0fbqvU6mi859D; reg [6:0] DOFNWCpbdQSLsWtzwny1qG; reg EWvO8Kf2QN2SS53GJJcWwF; reg [2:0] j9HNozHmNa6lYL8HVho1pB; reg B9qRWWVXUMKaf08lKjOj5G; wire signed [15:0] zVla2Vy8BUCugJ5Gig2ZK [0:127]; wire signed [15:0] F8NQxbAEqqIEtFo6mesHd; reg signed [15:0] CIRDDBHrGgCpm7HNrbXUCF; wire signed [15:0] ysWUViVY5R4DChvjvp5gDD [0:127]; wire signed [15:0] jsn1oqDToTuWwgUlIvqN3; reg signed [15:0] M9MMs7oRisnNmiBXjmtOsD; reg [2:0] YjlT6Mg9KMpPzxF47HzV7D; reg UrNpVdQvuAmKReKH4NECKD; reg signed [15:0] xiCPrrY7lS0ezOvEYWzkuG; reg signed [15:0] KlnKP5IsEqVnpuj6nZXNwC; reg [2:0] CbpoQEK97vFu56nv3223yC; reg [9:0] ZWvsxRFpFAzxN5xMmZuitE; reg signed [21:0] uCEkpKGKs7tQvr2GeEGSGC; reg signed [21:0] hhzTcPgpleSJBYLOoujKGG; reg signed [11:0] cVX5EXK4yxLZ1cYzNgyXx; reg signed [11:0] g4zMZYWhK020aMvVlufXSO; reg signed [21:0] SVYTAuHmM7AdeQD3dklB3D; reg signed [21:0] z9uPanlNUawhpWBfZzoV6C; reg signed [21:0] iKPA1JOFbNoLsuo87UbsvD; reg signed [21:0] K3fvtqFABfYnMEzDvYIrq; reg signed [11:0] jbCFxKpbanHjkeuxNFuv1D; reg signed [11:0] xs6NJDxbN0KSgBeqxxDWYF; reg signed [15:0] KwiyVhhhZdTrDQCbiLV8zE; reg signed [15:0] sGNGvuvL8Q7LZvZSVKC57B; reg signed [16:0] WJY0hyRMua5sU8DuMmLu4; reg signed [16:0] b6ofl8SS59auHuq7NOO0WOG; reg signed [16:0] f2RPd8CpcTyQnKsmtWEywG; reg signed [16:0] w4sUCJ8sn9dqukS5aRJDigE; reg signed [16:0] L3USkDc1T9xpZF6CkNG03D; reg signed [16:0] s195ulFHSeSTCYTLhumIdD; wire Yftze0y14b5d5HigFNuUBH; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : A7mAa8MkEw1SBVJbtTHnZE if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin URO3uEJ9VVi4n2rv5pG4XF <= 3'b000; mevVutOyAH9CPJEBvvvxsF <= 10'b0000000000; Mndh5cWFT2MK7irxEkUgvB <= 7'b0000000; DSwbuqNl6si2qBBlHlS4m <= 1'b0; ADYssd29ifP9Cnqtxk4KFH <= 1'b0; zUwvjmWVganUujWHX9Ik8G <= 1'b0; TE2s9kaW4jbT2yuidpcUIF <= 8'b00000000; j9GInQQXHbUGPAy0R0X4BQD <= 2'b00; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin URO3uEJ9VVi4n2rv5pG4XF <= 3'b000; mevVutOyAH9CPJEBvvvxsF <= 10'b0000000000; Mndh5cWFT2MK7irxEkUgvB <= 7'b0000000; DSwbuqNl6si2qBBlHlS4m <= 1'b0; ADYssd29ifP9Cnqtxk4KFH <= 1'b0; zUwvjmWVganUujWHX9Ik8G <= 1'b0; TE2s9kaW4jbT2yuidpcUIF <= 8'b00000000; j9GInQQXHbUGPAy0R0X4BQD <= 2'b00; end else begin TE2s9kaW4jbT2yuidpcUIF <= vyYw1SbJbcSwGlwsC50cRF; j9GInQQXHbUGPAy0R0X4BQD <= tHBJR87iWmyApKoUBwoC; URO3uEJ9VVi4n2rv5pG4XF <= ZXzEhgRyMkDiwOKQ1ZyHtH; mevVutOyAH9CPJEBvvvxsF <= vndcJtBZasetzBa7iOZamH; Mndh5cWFT2MK7irxEkUgvB <= W3LV4fQGt3vLDwUnzRRUwH; DSwbuqNl6si2qBBlHlS4m <= t96JNxh4AbzBXPo2zT29dlG; ADYssd29ifP9Cnqtxk4KFH <= ARo3kgZ8gBa9Exsckya1UB; zUwvjmWVganUujWHX9Ik8G <= IvvfGB2My0fbqvU6mi859D; end end end always @(ADYssd29ifP9Cnqtxk4KFH, DSwbuqNl6si2qBBlHlS4m, Mndh5cWFT2MK7irxEkUgvB, NMWfejbHi1tIjFkylFWDkC, TE2s9kaW4jbT2yuidpcUIF, URO3uEJ9VVi4n2rv5pG4XF, j9GInQQXHbUGPAy0R0X4BQD, mevVutOyAH9CPJEBvvvxsF, zUwvjmWVganUujWHX9Ik8G) begin hhzTcPgpleSJBYLOoujKGG = 22'sb0000000000000000000000; cVX5EXK4yxLZ1cYzNgyXx = 12'sb000000000000; g4zMZYWhK020aMvVlufXSO = 12'sb000000000000; z9uPanlNUawhpWBfZzoV6C = 22'sb0000000000000000000000; K3fvtqFABfYnMEzDvYIrq = 22'sb0000000000000000000000; ZWvsxRFpFAzxN5xMmZuitE = 10'b0000000000; uCEkpKGKs7tQvr2GeEGSGC = 22'sb0000000000000000000000; SVYTAuHmM7AdeQD3dklB3D = 22'sb0000000000000000000000; iKPA1JOFbNoLsuo87UbsvD = 22'sb0000000000000000000000; jbCFxKpbanHjkeuxNFuv1D = 12'sb000000000000; xs6NJDxbN0KSgBeqxxDWYF = 12'sb000000000000; vyYw1SbJbcSwGlwsC50cRF = TE2s9kaW4jbT2yuidpcUIF; tHBJR87iWmyApKoUBwoC = j9GInQQXHbUGPAy0R0X4BQD; vndcJtBZasetzBa7iOZamH = mevVutOyAH9CPJEBvvvxsF; W3LV4fQGt3vLDwUnzRRUwH = Mndh5cWFT2MK7irxEkUgvB; t96JNxh4AbzBXPo2zT29dlG = DSwbuqNl6si2qBBlHlS4m; IvvfGB2My0fbqvU6mi859D = ADYssd29ifP9Cnqtxk4KFH; ARo3kgZ8gBa9Exsckya1UB = NMWfejbHi1tIjFkylFWDkC; case ( mevVutOyAH9CPJEBvvvxsF) 10'b0010000000 : begin CbpoQEK97vFu56nv3223yC = 3'b000; t96JNxh4AbzBXPo2zT29dlG = 1'b1; end 10'b0100000000 : begin CbpoQEK97vFu56nv3223yC = 3'b001; t96JNxh4AbzBXPo2zT29dlG = 1'b0; end 10'b0110000000 : begin CbpoQEK97vFu56nv3223yC = 3'b010; t96JNxh4AbzBXPo2zT29dlG = 1'b1; end 10'b1000000000 : begin CbpoQEK97vFu56nv3223yC = 3'b011; t96JNxh4AbzBXPo2zT29dlG = 1'b0; end 10'b1010000000 : begin CbpoQEK97vFu56nv3223yC = 3'b100; t96JNxh4AbzBXPo2zT29dlG = 1'b1; end default : begin CbpoQEK97vFu56nv3223yC = mevVutOyAH9CPJEBvvvxsF[9:7]; t96JNxh4AbzBXPo2zT29dlG = 1'b0; end endcase ZXzEhgRyMkDiwOKQ1ZyHtH = CbpoQEK97vFu56nv3223yC; case ( CbpoQEK97vFu56nv3223yC) 3'b000 : begin W3LV4fQGt3vLDwUnzRRUwH = mevVutOyAH9CPJEBvvvxsF[6:0]; end 3'b001 : begin jbCFxKpbanHjkeuxNFuv1D = {2'b0, mevVutOyAH9CPJEBvvvxsF}; cVX5EXK4yxLZ1cYzNgyXx = 12'sb000100000000 - jbCFxKpbanHjkeuxNFuv1D; W3LV4fQGt3vLDwUnzRRUwH = cVX5EXK4yxLZ1cYzNgyXx[6:0]; end 3'b010 : begin xs6NJDxbN0KSgBeqxxDWYF = {2'b0, mevVutOyAH9CPJEBvvvxsF}; g4zMZYWhK020aMvVlufXSO = xs6NJDxbN0KSgBeqxxDWYF - 12'sb000100000000; W3LV4fQGt3vLDwUnzRRUwH = g4zMZYWhK020aMvVlufXSO[6:0]; end 3'b011 : begin SVYTAuHmM7AdeQD3dklB3D = {5'b0, {mevVutOyAH9CPJEBvvvxsF, 7'b0000000}}; z9uPanlNUawhpWBfZzoV6C = 22'sb0000010000000000000000 - SVYTAuHmM7AdeQD3dklB3D; W3LV4fQGt3vLDwUnzRRUwH = z9uPanlNUawhpWBfZzoV6C[13:7]; end 3'b100 : begin iKPA1JOFbNoLsuo87UbsvD = {5'b0, {mevVutOyAH9CPJEBvvvxsF, 7'b0000000}}; K3fvtqFABfYnMEzDvYIrq = iKPA1JOFbNoLsuo87UbsvD - 22'sb0000010000000000000000; W3LV4fQGt3vLDwUnzRRUwH = K3fvtqFABfYnMEzDvYIrq[13:7]; end default : begin uCEkpKGKs7tQvr2GeEGSGC = {5'b0, {mevVutOyAH9CPJEBvvvxsF, 7'b0000000}}; hhzTcPgpleSJBYLOoujKGG = 22'sb0000011000000000000000 - uCEkpKGKs7tQvr2GeEGSGC; W3LV4fQGt3vLDwUnzRRUwH = hhzTcPgpleSJBYLOoujKGG[13:7]; end endcase if (j9GInQQXHbUGPAy0R0X4BQD == 2'b00) begin vndcJtBZasetzBa7iOZamH = 10'b0000000000; end else if (j9GInQQXHbUGPAy0R0X4BQD == 2'b01) begin vndcJtBZasetzBa7iOZamH = {2'b0, TE2s9kaW4jbT2yuidpcUIF} <<< 8'd1; end else if (j9GInQQXHbUGPAy0R0X4BQD == 2'b10) begin vndcJtBZasetzBa7iOZamH = {2'b0, TE2s9kaW4jbT2yuidpcUIF}; end else begin ZWvsxRFpFAzxN5xMmZuitE = {2'b0, TE2s9kaW4jbT2yuidpcUIF}; vndcJtBZasetzBa7iOZamH = (ZWvsxRFpFAzxN5xMmZuitE <<< 8'd1) + ZWvsxRFpFAzxN5xMmZuitE; end if (NMWfejbHi1tIjFkylFWDkC && (TE2s9kaW4jbT2yuidpcUIF > 8'b11101111)) begin tHBJR87iWmyApKoUBwoC = j9GInQQXHbUGPAy0R0X4BQD + 2'b01; end if (NMWfejbHi1tIjFkylFWDkC) begin vyYw1SbJbcSwGlwsC50cRF = TE2s9kaW4jbT2yuidpcUIF + 8'b00010000; end DOFNWCpbdQSLsWtzwny1qG = Mndh5cWFT2MK7irxEkUgvB; EWvO8Kf2QN2SS53GJJcWwF = zUwvjmWVganUujWHX9Ik8G; j9HNozHmNa6lYL8HVho1pB = URO3uEJ9VVi4n2rv5pG4XF; B9qRWWVXUMKaf08lKjOj5G = DSwbuqNl6si2qBBlHlS4m; end assign zVla2Vy8BUCugJ5Gig2ZK[0] = 16'sb0100000000000000; assign zVla2Vy8BUCugJ5Gig2ZK[1] = 16'sb0100000000000000; assign zVla2Vy8BUCugJ5Gig2ZK[2] = 16'sb0011111111111111; assign zVla2Vy8BUCugJ5Gig2ZK[3] = 16'sb0011111111111101; assign zVla2Vy8BUCugJ5Gig2ZK[4] = 16'sb0011111111111011; assign zVla2Vy8BUCugJ5Gig2ZK[5] = 16'sb0011111111111000; assign zVla2Vy8BUCugJ5Gig2ZK[6] = 16'sb0011111111110101; assign zVla2Vy8BUCugJ5Gig2ZK[7] = 16'sb0011111111110001; assign zVla2Vy8BUCugJ5Gig2ZK[8] = 16'sb0011111111101100; assign zVla2Vy8BUCugJ5Gig2ZK[9] = 16'sb0011111111100111; assign zVla2Vy8BUCugJ5Gig2ZK[10] = 16'sb0011111111100001; assign zVla2Vy8BUCugJ5Gig2ZK[11] = 16'sb0011111111011011; assign zVla2Vy8BUCugJ5Gig2ZK[12] = 16'sb0011111111010100; assign zVla2Vy8BUCugJ5Gig2ZK[13] = 16'sb0011111111001100; assign zVla2Vy8BUCugJ5Gig2ZK[14] = 16'sb0011111111000100; assign zVla2Vy8BUCugJ5Gig2ZK[15] = 16'sb0011111110111011; assign zVla2Vy8BUCugJ5Gig2ZK[16] = 16'sb0011111110110001; assign zVla2Vy8BUCugJ5Gig2ZK[17] = 16'sb0011111110100111; assign zVla2Vy8BUCugJ5Gig2ZK[18] = 16'sb0011111110011100; assign zVla2Vy8BUCugJ5Gig2ZK[19] = 16'sb0011111110010001; assign zVla2Vy8BUCugJ5Gig2ZK[20] = 16'sb0011111110000101; assign zVla2Vy8BUCugJ5Gig2ZK[21] = 16'sb0011111101111000; assign zVla2Vy8BUCugJ5Gig2ZK[22] = 16'sb0011111101101011; assign zVla2Vy8BUCugJ5Gig2ZK[23] = 16'sb0011111101011101; assign zVla2Vy8BUCugJ5Gig2ZK[24] = 16'sb0011111101001111; assign zVla2Vy8BUCugJ5Gig2ZK[25] = 16'sb0011111101000000; assign zVla2Vy8BUCugJ5Gig2ZK[26] = 16'sb0011111100110000; assign zVla2Vy8BUCugJ5Gig2ZK[27] = 16'sb0011111100100000; assign zVla2Vy8BUCugJ5Gig2ZK[28] = 16'sb0011111100001111; assign zVla2Vy8BUCugJ5Gig2ZK[29] = 16'sb0011111011111101; assign zVla2Vy8BUCugJ5Gig2ZK[30] = 16'sb0011111011101011; assign zVla2Vy8BUCugJ5Gig2ZK[31] = 16'sb0011111011011000; assign zVla2Vy8BUCugJ5Gig2ZK[32] = 16'sb0011111011000101; assign zVla2Vy8BUCugJ5Gig2ZK[33] = 16'sb0011111010110001; assign zVla2Vy8BUCugJ5Gig2ZK[34] = 16'sb0011111010011101; assign zVla2Vy8BUCugJ5Gig2ZK[35] = 16'sb0011111010001000; assign zVla2Vy8BUCugJ5Gig2ZK[36] = 16'sb0011111001110010; assign zVla2Vy8BUCugJ5Gig2ZK[37] = 16'sb0011111001011100; assign zVla2Vy8BUCugJ5Gig2ZK[38] = 16'sb0011111001000101; assign zVla2Vy8BUCugJ5Gig2ZK[39] = 16'sb0011111000101101; assign zVla2Vy8BUCugJ5Gig2ZK[40] = 16'sb0011111000010101; assign zVla2Vy8BUCugJ5Gig2ZK[41] = 16'sb0011110111111100; assign zVla2Vy8BUCugJ5Gig2ZK[42] = 16'sb0011110111100011; assign zVla2Vy8BUCugJ5Gig2ZK[43] = 16'sb0011110111001001; assign zVla2Vy8BUCugJ5Gig2ZK[44] = 16'sb0011110110101111; assign zVla2Vy8BUCugJ5Gig2ZK[45] = 16'sb0011110110010011; assign zVla2Vy8BUCugJ5Gig2ZK[46] = 16'sb0011110101111000; assign zVla2Vy8BUCugJ5Gig2ZK[47] = 16'sb0011110101011011; assign zVla2Vy8BUCugJ5Gig2ZK[48] = 16'sb0011110100111111; assign zVla2Vy8BUCugJ5Gig2ZK[49] = 16'sb0011110100100001; assign zVla2Vy8BUCugJ5Gig2ZK[50] = 16'sb0011110100000011; assign zVla2Vy8BUCugJ5Gig2ZK[51] = 16'sb0011110011100100; assign zVla2Vy8BUCugJ5Gig2ZK[52] = 16'sb0011110011000101; assign zVla2Vy8BUCugJ5Gig2ZK[53] = 16'sb0011110010100101; assign zVla2Vy8BUCugJ5Gig2ZK[54] = 16'sb0011110010000101; assign zVla2Vy8BUCugJ5Gig2ZK[55] = 16'sb0011110001100100; assign zVla2Vy8BUCugJ5Gig2ZK[56] = 16'sb0011110001000010; assign zVla2Vy8BUCugJ5Gig2ZK[57] = 16'sb0011110000100000; assign zVla2Vy8BUCugJ5Gig2ZK[58] = 16'sb0011101111111101; assign zVla2Vy8BUCugJ5Gig2ZK[59] = 16'sb0011101111011010; assign zVla2Vy8BUCugJ5Gig2ZK[60] = 16'sb0011101110110110; assign zVla2Vy8BUCugJ5Gig2ZK[61] = 16'sb0011101110010010; assign zVla2Vy8BUCugJ5Gig2ZK[62] = 16'sb0011101101101101; assign zVla2Vy8BUCugJ5Gig2ZK[63] = 16'sb0011101101000111; assign zVla2Vy8BUCugJ5Gig2ZK[64] = 16'sb0011101100100001; assign zVla2Vy8BUCugJ5Gig2ZK[65] = 16'sb0011101011111010; assign zVla2Vy8BUCugJ5Gig2ZK[66] = 16'sb0011101011010011; assign zVla2Vy8BUCugJ5Gig2ZK[67] = 16'sb0011101010101011; assign zVla2Vy8BUCugJ5Gig2ZK[68] = 16'sb0011101010000010; assign zVla2Vy8BUCugJ5Gig2ZK[69] = 16'sb0011101001011001; assign zVla2Vy8BUCugJ5Gig2ZK[70] = 16'sb0011101000110000; assign zVla2Vy8BUCugJ5Gig2ZK[71] = 16'sb0011101000000110; assign zVla2Vy8BUCugJ5Gig2ZK[72] = 16'sb0011100111011011; assign zVla2Vy8BUCugJ5Gig2ZK[73] = 16'sb0011100110110000; assign zVla2Vy8BUCugJ5Gig2ZK[74] = 16'sb0011100110000100; assign zVla2Vy8BUCugJ5Gig2ZK[75] = 16'sb0011100101011000; assign zVla2Vy8BUCugJ5Gig2ZK[76] = 16'sb0011100100101011; assign zVla2Vy8BUCugJ5Gig2ZK[77] = 16'sb0011100011111101; assign zVla2Vy8BUCugJ5Gig2ZK[78] = 16'sb0011100011001111; assign zVla2Vy8BUCugJ5Gig2ZK[79] = 16'sb0011100010100001; assign zVla2Vy8BUCugJ5Gig2ZK[80] = 16'sb0011100001110001; assign zVla2Vy8BUCugJ5Gig2ZK[81] = 16'sb0011100001000010; assign zVla2Vy8BUCugJ5Gig2ZK[82] = 16'sb0011100000010010; assign zVla2Vy8BUCugJ5Gig2ZK[83] = 16'sb0011011111100001; assign zVla2Vy8BUCugJ5Gig2ZK[84] = 16'sb0011011110110000; assign zVla2Vy8BUCugJ5Gig2ZK[85] = 16'sb0011011101111110; assign zVla2Vy8BUCugJ5Gig2ZK[86] = 16'sb0011011101001011; assign zVla2Vy8BUCugJ5Gig2ZK[87] = 16'sb0011011100011000; assign zVla2Vy8BUCugJ5Gig2ZK[88] = 16'sb0011011011100101; assign zVla2Vy8BUCugJ5Gig2ZK[89] = 16'sb0011011010110001; assign zVla2Vy8BUCugJ5Gig2ZK[90] = 16'sb0011011001111101; assign zVla2Vy8BUCugJ5Gig2ZK[91] = 16'sb0011011001001000; assign zVla2Vy8BUCugJ5Gig2ZK[92] = 16'sb0011011000010010; assign zVla2Vy8BUCugJ5Gig2ZK[93] = 16'sb0011010111011100; assign zVla2Vy8BUCugJ5Gig2ZK[94] = 16'sb0011010110100101; assign zVla2Vy8BUCugJ5Gig2ZK[95] = 16'sb0011010101101110; assign zVla2Vy8BUCugJ5Gig2ZK[96] = 16'sb0011010100110111; assign zVla2Vy8BUCugJ5Gig2ZK[97] = 16'sb0011010011111111; assign zVla2Vy8BUCugJ5Gig2ZK[98] = 16'sb0011010011000110; assign zVla2Vy8BUCugJ5Gig2ZK[99] = 16'sb0011010010001101; assign zVla2Vy8BUCugJ5Gig2ZK[100] = 16'sb0011010001010011; assign zVla2Vy8BUCugJ5Gig2ZK[101] = 16'sb0011010000011001; assign zVla2Vy8BUCugJ5Gig2ZK[102] = 16'sb0011001111011111; assign zVla2Vy8BUCugJ5Gig2ZK[103] = 16'sb0011001110100011; assign zVla2Vy8BUCugJ5Gig2ZK[104] = 16'sb0011001101101000; assign zVla2Vy8BUCugJ5Gig2ZK[105] = 16'sb0011001100101100; assign zVla2Vy8BUCugJ5Gig2ZK[106] = 16'sb0011001011101111; assign zVla2Vy8BUCugJ5Gig2ZK[107] = 16'sb0011001010110010; assign zVla2Vy8BUCugJ5Gig2ZK[108] = 16'sb0011001001110100; assign zVla2Vy8BUCugJ5Gig2ZK[109] = 16'sb0011001000110110; assign zVla2Vy8BUCugJ5Gig2ZK[110] = 16'sb0011000111111000; assign zVla2Vy8BUCugJ5Gig2ZK[111] = 16'sb0011000110111001; assign zVla2Vy8BUCugJ5Gig2ZK[112] = 16'sb0011000101111001; assign zVla2Vy8BUCugJ5Gig2ZK[113] = 16'sb0011000100111001; assign zVla2Vy8BUCugJ5Gig2ZK[114] = 16'sb0011000011111001; assign zVla2Vy8BUCugJ5Gig2ZK[115] = 16'sb0011000010111000; assign zVla2Vy8BUCugJ5Gig2ZK[116] = 16'sb0011000001110110; assign zVla2Vy8BUCugJ5Gig2ZK[117] = 16'sb0011000000110100; assign zVla2Vy8BUCugJ5Gig2ZK[118] = 16'sb0010111111110010; assign zVla2Vy8BUCugJ5Gig2ZK[119] = 16'sb0010111110101111; assign zVla2Vy8BUCugJ5Gig2ZK[120] = 16'sb0010111101101100; assign zVla2Vy8BUCugJ5Gig2ZK[121] = 16'sb0010111100101000; assign zVla2Vy8BUCugJ5Gig2ZK[122] = 16'sb0010111011100100; assign zVla2Vy8BUCugJ5Gig2ZK[123] = 16'sb0010111010011111; assign zVla2Vy8BUCugJ5Gig2ZK[124] = 16'sb0010111001011010; assign zVla2Vy8BUCugJ5Gig2ZK[125] = 16'sb0010111000010101; assign zVla2Vy8BUCugJ5Gig2ZK[126] = 16'sb0010110111001111; assign zVla2Vy8BUCugJ5Gig2ZK[127] = 16'sb0010110110001000; assign F8NQxbAEqqIEtFo6mesHd = zVla2Vy8BUCugJ5Gig2ZK[DOFNWCpbdQSLsWtzwny1qG]; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : j0boDGRQkCezKyDxbtKinG if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin CIRDDBHrGgCpm7HNrbXUCF <= 16'sb0000000000000000; end else begin CIRDDBHrGgCpm7HNrbXUCF <= F8NQxbAEqqIEtFo6mesHd; end end assign ysWUViVY5R4DChvjvp5gDD[0] = 16'sb0000000000000000; assign ysWUViVY5R4DChvjvp5gDD[1] = 16'sb1111111110011011; assign ysWUViVY5R4DChvjvp5gDD[2] = 16'sb1111111100110111; assign ysWUViVY5R4DChvjvp5gDD[3] = 16'sb1111111011010010; assign ysWUViVY5R4DChvjvp5gDD[4] = 16'sb1111111001101110; assign ysWUViVY5R4DChvjvp5gDD[5] = 16'sb1111111000001001; assign ysWUViVY5R4DChvjvp5gDD[6] = 16'sb1111110110100101; assign ysWUViVY5R4DChvjvp5gDD[7] = 16'sb1111110101000000; assign ysWUViVY5R4DChvjvp5gDD[8] = 16'sb1111110011011100; assign ysWUViVY5R4DChvjvp5gDD[9] = 16'sb1111110001111000; assign ysWUViVY5R4DChvjvp5gDD[10] = 16'sb1111110000010011; assign ysWUViVY5R4DChvjvp5gDD[11] = 16'sb1111101110101111; assign ysWUViVY5R4DChvjvp5gDD[12] = 16'sb1111101101001011; assign ysWUViVY5R4DChvjvp5gDD[13] = 16'sb1111101011100110; assign ysWUViVY5R4DChvjvp5gDD[14] = 16'sb1111101010000010; assign ysWUViVY5R4DChvjvp5gDD[15] = 16'sb1111101000011110; assign ysWUViVY5R4DChvjvp5gDD[16] = 16'sb1111100110111010; assign ysWUViVY5R4DChvjvp5gDD[17] = 16'sb1111100101010110; assign ysWUViVY5R4DChvjvp5gDD[18] = 16'sb1111100011110010; assign ysWUViVY5R4DChvjvp5gDD[19] = 16'sb1111100010001110; assign ysWUViVY5R4DChvjvp5gDD[20] = 16'sb1111100000101010; assign ysWUViVY5R4DChvjvp5gDD[21] = 16'sb1111011111000111; assign ysWUViVY5R4DChvjvp5gDD[22] = 16'sb1111011101100011; assign ysWUViVY5R4DChvjvp5gDD[23] = 16'sb1111011011111111; assign ysWUViVY5R4DChvjvp5gDD[24] = 16'sb1111011010011100; assign ysWUViVY5R4DChvjvp5gDD[25] = 16'sb1111011000111001; assign ysWUViVY5R4DChvjvp5gDD[26] = 16'sb1111010111010101; assign ysWUViVY5R4DChvjvp5gDD[27] = 16'sb1111010101110010; assign ysWUViVY5R4DChvjvp5gDD[28] = 16'sb1111010100001111; assign ysWUViVY5R4DChvjvp5gDD[29] = 16'sb1111010010101100; assign ysWUViVY5R4DChvjvp5gDD[30] = 16'sb1111010001001001; assign ysWUViVY5R4DChvjvp5gDD[31] = 16'sb1111001111100110; assign ysWUViVY5R4DChvjvp5gDD[32] = 16'sb1111001110000100; assign ysWUViVY5R4DChvjvp5gDD[33] = 16'sb1111001100100001; assign ysWUViVY5R4DChvjvp5gDD[34] = 16'sb1111001010111111; assign ysWUViVY5R4DChvjvp5gDD[35] = 16'sb1111001001011100; assign ysWUViVY5R4DChvjvp5gDD[36] = 16'sb1111000111111010; assign ysWUViVY5R4DChvjvp5gDD[37] = 16'sb1111000110011000; assign ysWUViVY5R4DChvjvp5gDD[38] = 16'sb1111000100110110; assign ysWUViVY5R4DChvjvp5gDD[39] = 16'sb1111000011010101; assign ysWUViVY5R4DChvjvp5gDD[40] = 16'sb1111000001110011; assign ysWUViVY5R4DChvjvp5gDD[41] = 16'sb1111000000010010; assign ysWUViVY5R4DChvjvp5gDD[42] = 16'sb1110111110110000; assign ysWUViVY5R4DChvjvp5gDD[43] = 16'sb1110111101001111; assign ysWUViVY5R4DChvjvp5gDD[44] = 16'sb1110111011101110; assign ysWUViVY5R4DChvjvp5gDD[45] = 16'sb1110111010001101; assign ysWUViVY5R4DChvjvp5gDD[46] = 16'sb1110111000101101; assign ysWUViVY5R4DChvjvp5gDD[47] = 16'sb1110110111001100; assign ysWUViVY5R4DChvjvp5gDD[48] = 16'sb1110110101101100; assign ysWUViVY5R4DChvjvp5gDD[49] = 16'sb1110110100001100; assign ysWUViVY5R4DChvjvp5gDD[50] = 16'sb1110110010101100; assign ysWUViVY5R4DChvjvp5gDD[51] = 16'sb1110110001001100; assign ysWUViVY5R4DChvjvp5gDD[52] = 16'sb1110101111101101; assign ysWUViVY5R4DChvjvp5gDD[53] = 16'sb1110101110001101; assign ysWUViVY5R4DChvjvp5gDD[54] = 16'sb1110101100101110; assign ysWUViVY5R4DChvjvp5gDD[55] = 16'sb1110101011001111; assign ysWUViVY5R4DChvjvp5gDD[56] = 16'sb1110101001110000; assign ysWUViVY5R4DChvjvp5gDD[57] = 16'sb1110101000010010; assign ysWUViVY5R4DChvjvp5gDD[58] = 16'sb1110100110110100; assign ysWUViVY5R4DChvjvp5gDD[59] = 16'sb1110100101010101; assign ysWUViVY5R4DChvjvp5gDD[60] = 16'sb1110100011110111; assign ysWUViVY5R4DChvjvp5gDD[61] = 16'sb1110100010011010; assign ysWUViVY5R4DChvjvp5gDD[62] = 16'sb1110100000111100; assign ysWUViVY5R4DChvjvp5gDD[63] = 16'sb1110011111011111; assign ysWUViVY5R4DChvjvp5gDD[64] = 16'sb1110011110000010; assign ysWUViVY5R4DChvjvp5gDD[65] = 16'sb1110011100100101; assign ysWUViVY5R4DChvjvp5gDD[66] = 16'sb1110011011001001; assign ysWUViVY5R4DChvjvp5gDD[67] = 16'sb1110011001101101; assign ysWUViVY5R4DChvjvp5gDD[68] = 16'sb1110011000010001; assign ysWUViVY5R4DChvjvp5gDD[69] = 16'sb1110010110110101; assign ysWUViVY5R4DChvjvp5gDD[70] = 16'sb1110010101011001; assign ysWUViVY5R4DChvjvp5gDD[71] = 16'sb1110010011111110; assign ysWUViVY5R4DChvjvp5gDD[72] = 16'sb1110010010100011; assign ysWUViVY5R4DChvjvp5gDD[73] = 16'sb1110010001001000; assign ysWUViVY5R4DChvjvp5gDD[74] = 16'sb1110001111101110; assign ysWUViVY5R4DChvjvp5gDD[75] = 16'sb1110001110010100; assign ysWUViVY5R4DChvjvp5gDD[76] = 16'sb1110001100111010; assign ysWUViVY5R4DChvjvp5gDD[77] = 16'sb1110001011100000; assign ysWUViVY5R4DChvjvp5gDD[78] = 16'sb1110001010000111; assign ysWUViVY5R4DChvjvp5gDD[79] = 16'sb1110001000101101; assign ysWUViVY5R4DChvjvp5gDD[80] = 16'sb1110000111010101; assign ysWUViVY5R4DChvjvp5gDD[81] = 16'sb1110000101111100; assign ysWUViVY5R4DChvjvp5gDD[82] = 16'sb1110000100100100; assign ysWUViVY5R4DChvjvp5gDD[83] = 16'sb1110000011001100; assign ysWUViVY5R4DChvjvp5gDD[84] = 16'sb1110000001110100; assign ysWUViVY5R4DChvjvp5gDD[85] = 16'sb1110000000011101; assign ysWUViVY5R4DChvjvp5gDD[86] = 16'sb1101111111000110; assign ysWUViVY5R4DChvjvp5gDD[87] = 16'sb1101111101101111; assign ysWUViVY5R4DChvjvp5gDD[88] = 16'sb1101111100011001; assign ysWUViVY5R4DChvjvp5gDD[89] = 16'sb1101111011000011; assign ysWUViVY5R4DChvjvp5gDD[90] = 16'sb1101111001101101; assign ysWUViVY5R4DChvjvp5gDD[91] = 16'sb1101111000011000; assign ysWUViVY5R4DChvjvp5gDD[92] = 16'sb1101110111000011; assign ysWUViVY5R4DChvjvp5gDD[93] = 16'sb1101110101101110; assign ysWUViVY5R4DChvjvp5gDD[94] = 16'sb1101110100011001; assign ysWUViVY5R4DChvjvp5gDD[95] = 16'sb1101110011000101; assign ysWUViVY5R4DChvjvp5gDD[96] = 16'sb1101110001110010; assign ysWUViVY5R4DChvjvp5gDD[97] = 16'sb1101110000011110; assign ysWUViVY5R4DChvjvp5gDD[98] = 16'sb1101101111001011; assign ysWUViVY5R4DChvjvp5gDD[99] = 16'sb1101101101111000; assign ysWUViVY5R4DChvjvp5gDD[100] = 16'sb1101101100100110; assign ysWUViVY5R4DChvjvp5gDD[101] = 16'sb1101101011010100; assign ysWUViVY5R4DChvjvp5gDD[102] = 16'sb1101101010000010; assign ysWUViVY5R4DChvjvp5gDD[103] = 16'sb1101101000110001; assign ysWUViVY5R4DChvjvp5gDD[104] = 16'sb1101100111100000; assign ysWUViVY5R4DChvjvp5gDD[105] = 16'sb1101100110001111; assign ysWUViVY5R4DChvjvp5gDD[106] = 16'sb1101100100111111; assign ysWUViVY5R4DChvjvp5gDD[107] = 16'sb1101100011101111; assign ysWUViVY5R4DChvjvp5gDD[108] = 16'sb1101100010100000; assign ysWUViVY5R4DChvjvp5gDD[109] = 16'sb1101100001010001; assign ysWUViVY5R4DChvjvp5gDD[110] = 16'sb1101100000000010; assign ysWUViVY5R4DChvjvp5gDD[111] = 16'sb1101011110110100; assign ysWUViVY5R4DChvjvp5gDD[112] = 16'sb1101011101100110; assign ysWUViVY5R4DChvjvp5gDD[113] = 16'sb1101011100011001; assign ysWUViVY5R4DChvjvp5gDD[114] = 16'sb1101011011001011; assign ysWUViVY5R4DChvjvp5gDD[115] = 16'sb1101011001111111; assign ysWUViVY5R4DChvjvp5gDD[116] = 16'sb1101011000110010; assign ysWUViVY5R4DChvjvp5gDD[117] = 16'sb1101010111100110; assign ysWUViVY5R4DChvjvp5gDD[118] = 16'sb1101010110011011; assign ysWUViVY5R4DChvjvp5gDD[119] = 16'sb1101010101010000; assign ysWUViVY5R4DChvjvp5gDD[120] = 16'sb1101010100000101; assign ysWUViVY5R4DChvjvp5gDD[121] = 16'sb1101010010111011; assign ysWUViVY5R4DChvjvp5gDD[122] = 16'sb1101010001110001; assign ysWUViVY5R4DChvjvp5gDD[123] = 16'sb1101010000101000; assign ysWUViVY5R4DChvjvp5gDD[124] = 16'sb1101001111011111; assign ysWUViVY5R4DChvjvp5gDD[125] = 16'sb1101001110010110; assign ysWUViVY5R4DChvjvp5gDD[126] = 16'sb1101001101001110; assign ysWUViVY5R4DChvjvp5gDD[127] = 16'sb1101001100000110; assign jsn1oqDToTuWwgUlIvqN3 = ysWUViVY5R4DChvjvp5gDD[DOFNWCpbdQSLsWtzwny1qG]; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : VAVA4twBRLX2WfwOrbR5l if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin M9MMs7oRisnNmiBXjmtOsD <= 16'sb0000000000000000; end else begin M9MMs7oRisnNmiBXjmtOsD <= jsn1oqDToTuWwgUlIvqN3; end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : MczQYJ6MT1pYZD7C1UhQv if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin YjlT6Mg9KMpPzxF47HzV7D <= 3'b000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin YjlT6Mg9KMpPzxF47HzV7D <= 3'b000; end else begin YjlT6Mg9KMpPzxF47HzV7D <= j9HNozHmNa6lYL8HVho1pB; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : xwyxj2YIc64Lxvl4r8S8mG if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin UrNpVdQvuAmKReKH4NECKD <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin UrNpVdQvuAmKReKH4NECKD <= 1'b0; end else begin UrNpVdQvuAmKReKH4NECKD <= B9qRWWVXUMKaf08lKjOj5G; end end end always @(CIRDDBHrGgCpm7HNrbXUCF, M9MMs7oRisnNmiBXjmtOsD, UrNpVdQvuAmKReKH4NECKD, YjlT6Mg9KMpPzxF47HzV7D) begin WJY0hyRMua5sU8DuMmLu4 = 17'sb00000000000000000; b6ofl8SS59auHuq7NOO0WOG = 17'sb00000000000000000; f2RPd8CpcTyQnKsmtWEywG = 17'sb00000000000000000; w4sUCJ8sn9dqukS5aRJDigE = 17'sb00000000000000000; L3USkDc1T9xpZF6CkNG03D = 17'sb00000000000000000; s195ulFHSeSTCYTLhumIdD = 17'sb00000000000000000; KwiyVhhhZdTrDQCbiLV8zE = CIRDDBHrGgCpm7HNrbXUCF; sGNGvuvL8Q7LZvZSVKC57B = M9MMs7oRisnNmiBXjmtOsD; if (UrNpVdQvuAmKReKH4NECKD) begin case ( YjlT6Mg9KMpPzxF47HzV7D) 3'b000 : begin KwiyVhhhZdTrDQCbiLV8zE = 16'sb0010110101000001; sGNGvuvL8Q7LZvZSVKC57B = 16'sb1101001010111111; end 3'b010 : begin KwiyVhhhZdTrDQCbiLV8zE = 16'sb1101001010111111; sGNGvuvL8Q7LZvZSVKC57B = 16'sb1101001010111111; end 3'b100 : begin KwiyVhhhZdTrDQCbiLV8zE = 16'sb1101001010111111; sGNGvuvL8Q7LZvZSVKC57B = 16'sb0010110101000001; end default : begin KwiyVhhhZdTrDQCbiLV8zE = 16'sb0010110101000001; sGNGvuvL8Q7LZvZSVKC57B = 16'sb1101001010111111; end endcase end else begin case ( YjlT6Mg9KMpPzxF47HzV7D) 3'b000 : begin end 3'b001 : begin WJY0hyRMua5sU8DuMmLu4 = - ({M9MMs7oRisnNmiBXjmtOsD[15], M9MMs7oRisnNmiBXjmtOsD}); KwiyVhhhZdTrDQCbiLV8zE = WJY0hyRMua5sU8DuMmLu4[15:0]; w4sUCJ8sn9dqukS5aRJDigE = - ({CIRDDBHrGgCpm7HNrbXUCF[15], CIRDDBHrGgCpm7HNrbXUCF}); sGNGvuvL8Q7LZvZSVKC57B = w4sUCJ8sn9dqukS5aRJDigE[15:0]; end 3'b010 : begin KwiyVhhhZdTrDQCbiLV8zE = M9MMs7oRisnNmiBXjmtOsD; L3USkDc1T9xpZF6CkNG03D = - ({CIRDDBHrGgCpm7HNrbXUCF[15], CIRDDBHrGgCpm7HNrbXUCF}); sGNGvuvL8Q7LZvZSVKC57B = L3USkDc1T9xpZF6CkNG03D[15:0]; end 3'b011 : begin b6ofl8SS59auHuq7NOO0WOG = - ({CIRDDBHrGgCpm7HNrbXUCF[15], CIRDDBHrGgCpm7HNrbXUCF}); KwiyVhhhZdTrDQCbiLV8zE = b6ofl8SS59auHuq7NOO0WOG[15:0]; sGNGvuvL8Q7LZvZSVKC57B = M9MMs7oRisnNmiBXjmtOsD; end 3'b100 : begin f2RPd8CpcTyQnKsmtWEywG = - ({CIRDDBHrGgCpm7HNrbXUCF[15], CIRDDBHrGgCpm7HNrbXUCF}); KwiyVhhhZdTrDQCbiLV8zE = f2RPd8CpcTyQnKsmtWEywG[15:0]; s195ulFHSeSTCYTLhumIdD = - ({M9MMs7oRisnNmiBXjmtOsD[15], M9MMs7oRisnNmiBXjmtOsD}); sGNGvuvL8Q7LZvZSVKC57B = s195ulFHSeSTCYTLhumIdD[15:0]; end default : begin KwiyVhhhZdTrDQCbiLV8zE = M9MMs7oRisnNmiBXjmtOsD; sGNGvuvL8Q7LZvZSVKC57B = CIRDDBHrGgCpm7HNrbXUCF; end endcase end xiCPrrY7lS0ezOvEYWzkuG = KwiyVhhhZdTrDQCbiLV8zE; KlnKP5IsEqVnpuj6nZXNwC = sGNGvuvL8Q7LZvZSVKC57B; end assign HXT3YNFExOHI94Xq9VVUBG = xiCPrrY7lS0ezOvEYWzkuG; assign EI1r2DTkmcgS5siR9DUFpG = KlnKP5IsEqVnpuj6nZXNwC; endmodule