`timescale 1 ns / 1 ns module CcegpoX8iivyKlrAI1PDCD (v04pHKxyc2sPW047bbyUgE, JAMOfrNHxGSYDF0urqkLN, EnlAo7K66kKuzHIKWLmc1F, ew3EeLap6s8rXmNrsqaTWH, qmhLAZZAHFrO09l1zXnPRC, JMtgCMT5TVzyJSn9uILA1, Z7ZDy0EvwvoCh1zahAqvSF, R6zf5iqRNVEGVBO8egq8kF, B58twvtfgVWGK5P29KavtH, qhk6Uhwhppvpssqm7Nh6XE, k3VfrgkD6DWITJL9WW5W4D, pPn6MVGqBLqJ0xzN2WYfFG, jNZ4xylBKAANfCL11XNxzB); input v04pHKxyc2sPW047bbyUgE; input JAMOfrNHxGSYDF0urqkLN; input signed [15:0] EnlAo7K66kKuzHIKWLmc1F; input signed [15:0] ew3EeLap6s8rXmNrsqaTWH; input signed [15:0] qmhLAZZAHFrO09l1zXnPRC; input signed [15:0] JMtgCMT5TVzyJSn9uILA1; input Z7ZDy0EvwvoCh1zahAqvSF; input R6zf5iqRNVEGVBO8egq8kF; output signed [15:0] B58twvtfgVWGK5P29KavtH; output signed [15:0] qhk6Uhwhppvpssqm7Nh6XE; output signed [15:0] k3VfrgkD6DWITJL9WW5W4D; output signed [15:0] pPn6MVGqBLqJ0xzN2WYfFG; output jNZ4xylBKAANfCL11XNxzB; reg signed [16:0] JuEdAzP84rg2g9z7jUH4CD; reg signed [16:0] w13lDdnHeKbz12RPLclXaYB; reg signed [16:0] G1cI3X0rnsuzwQl9n17YG; reg signed [16:0] GXg6LN8xFsDjdENYEDgKvC; reg c4yitNmVtLmJQVcYGJPLIKF; reg signed [16:0] EwpgnQRNtLL4vjPMlLBwS; reg signed [16:0] wf6CdozoYkNBecSlGbH3aH; reg signed [16:0] EVnidbw743875wavOVIR7C; reg signed [16:0] o238XHbXd6S5MNKr5zezYE; reg u3HkQauhqeq4XUajUjEhKC; reg signed [15:0] A5SQIaNgqW7DcTqQkKRVeD; reg signed [15:0] GaetbCaMty7UkzjqNoYErC; reg signed [15:0] M5AqS9R7rFTkWxwo8io2rH; reg signed [15:0] lcJo4MnEaj41ofRAtLkn4D; reg xijMuK2nBHoByB8rlrH50E; reg signed [16:0] sePOIYBEAAbt3DPar8jd5F; reg signed [16:0] iR0ShkyVRkHalUKTDnP0tG; reg signed [16:0] j3ureEigNPclVAPr6VwHVbG; reg signed [16:0] PmhJP7JCYGM2OStQXGIHgD; reg signed [16:0] TqfF3Zgxtm2cKWvwqij3m; reg signed [16:0] xijHKILnnZ8AgezrLRQvfF; reg signed [16:0] LoYaOvLnEQPAYlYtjywSTF; reg signed [16:0] Wf2SXd0xW1vBpZ49DhpQPE; reg signed [16:0] q5X9uuOdY7IBIroLr9svCOD; reg signed [16:0] BWK9w55Ml1WM8fecaddoXH; reg signed [16:0] h5B5oTxicZ5M23LhruZny; reg signed [16:0] DZuRxUKTwIbTxoU1h9ItHG; reg signed [16:0] pePHH82YpiwDZXNTNuW0kE; reg signed [16:0] w2JsFHlps9UnWS2sz8ntdrD; reg signed [16:0] Tyt8bZLXYY8su2Ax3b0rDH; reg signed [16:0] FZwXLiG4fwR5D6OFWbauRD; reg signed [16:0] b9TGb0JMaIybP28lLxuqbSD; reg signed [16:0] soGohDPw7ZeleH1CUwdFeD; reg signed [16:0] B8FsciuTU1IBtwPIKxFjdD; reg signed [16:0] V38Q9K9It91xb35KJJQllB; wire KTO4LzMG29up08DYwA89LE; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : cByCCMbEZEcgRtZNjjMl3D if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin JuEdAzP84rg2g9z7jUH4CD <= 17'sb00000000000000000; w13lDdnHeKbz12RPLclXaYB <= 17'sb00000000000000000; G1cI3X0rnsuzwQl9n17YG <= 17'sb00000000000000000; GXg6LN8xFsDjdENYEDgKvC <= 17'sb00000000000000000; c4yitNmVtLmJQVcYGJPLIKF <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin JuEdAzP84rg2g9z7jUH4CD <= 17'sb00000000000000000; w13lDdnHeKbz12RPLclXaYB <= 17'sb00000000000000000; G1cI3X0rnsuzwQl9n17YG <= 17'sb00000000000000000; GXg6LN8xFsDjdENYEDgKvC <= 17'sb00000000000000000; c4yitNmVtLmJQVcYGJPLIKF <= 1'b0; end else begin JuEdAzP84rg2g9z7jUH4CD <= EwpgnQRNtLL4vjPMlLBwS; w13lDdnHeKbz12RPLclXaYB <= wf6CdozoYkNBecSlGbH3aH; G1cI3X0rnsuzwQl9n17YG <= EVnidbw743875wavOVIR7C; GXg6LN8xFsDjdENYEDgKvC <= o238XHbXd6S5MNKr5zezYE; c4yitNmVtLmJQVcYGJPLIKF <= u3HkQauhqeq4XUajUjEhKC; end end end always @(EnlAo7K66kKuzHIKWLmc1F, G1cI3X0rnsuzwQl9n17YG, GXg6LN8xFsDjdENYEDgKvC, JMtgCMT5TVzyJSn9uILA1, JuEdAzP84rg2g9z7jUH4CD, Z7ZDy0EvwvoCh1zahAqvSF, c4yitNmVtLmJQVcYGJPLIKF, ew3EeLap6s8rXmNrsqaTWH, qmhLAZZAHFrO09l1zXnPRC, w13lDdnHeKbz12RPLclXaYB) begin pePHH82YpiwDZXNTNuW0kE = 17'sb00000000000000000; w2JsFHlps9UnWS2sz8ntdrD = 17'sb00000000000000000; Tyt8bZLXYY8su2Ax3b0rDH = 17'sb00000000000000000; FZwXLiG4fwR5D6OFWbauRD = 17'sb00000000000000000; b9TGb0JMaIybP28lLxuqbSD = 17'sb00000000000000000; soGohDPw7ZeleH1CUwdFeD = 17'sb00000000000000000; B8FsciuTU1IBtwPIKxFjdD = 17'sb00000000000000000; V38Q9K9It91xb35KJJQllB = 17'sb00000000000000000; EwpgnQRNtLL4vjPMlLBwS = JuEdAzP84rg2g9z7jUH4CD; wf6CdozoYkNBecSlGbH3aH = w13lDdnHeKbz12RPLclXaYB; EVnidbw743875wavOVIR7C = G1cI3X0rnsuzwQl9n17YG; o238XHbXd6S5MNKr5zezYE = GXg6LN8xFsDjdENYEDgKvC; u3HkQauhqeq4XUajUjEhKC = Z7ZDy0EvwvoCh1zahAqvSF; if (Z7ZDy0EvwvoCh1zahAqvSF) begin pePHH82YpiwDZXNTNuW0kE = {EnlAo7K66kKuzHIKWLmc1F[15], EnlAo7K66kKuzHIKWLmc1F}; w2JsFHlps9UnWS2sz8ntdrD = {qmhLAZZAHFrO09l1zXnPRC[15], qmhLAZZAHFrO09l1zXnPRC}; EwpgnQRNtLL4vjPMlLBwS = pePHH82YpiwDZXNTNuW0kE + w2JsFHlps9UnWS2sz8ntdrD; Tyt8bZLXYY8su2Ax3b0rDH = {EnlAo7K66kKuzHIKWLmc1F[15], EnlAo7K66kKuzHIKWLmc1F}; FZwXLiG4fwR5D6OFWbauRD = {qmhLAZZAHFrO09l1zXnPRC[15], qmhLAZZAHFrO09l1zXnPRC}; EVnidbw743875wavOVIR7C = Tyt8bZLXYY8su2Ax3b0rDH - FZwXLiG4fwR5D6OFWbauRD; b9TGb0JMaIybP28lLxuqbSD = {ew3EeLap6s8rXmNrsqaTWH[15], ew3EeLap6s8rXmNrsqaTWH}; soGohDPw7ZeleH1CUwdFeD = {JMtgCMT5TVzyJSn9uILA1[15], JMtgCMT5TVzyJSn9uILA1}; wf6CdozoYkNBecSlGbH3aH = b9TGb0JMaIybP28lLxuqbSD + soGohDPw7ZeleH1CUwdFeD; B8FsciuTU1IBtwPIKxFjdD = {ew3EeLap6s8rXmNrsqaTWH[15], ew3EeLap6s8rXmNrsqaTWH}; V38Q9K9It91xb35KJJQllB = {JMtgCMT5TVzyJSn9uILA1[15], JMtgCMT5TVzyJSn9uILA1}; o238XHbXd6S5MNKr5zezYE = B8FsciuTU1IBtwPIKxFjdD - V38Q9K9It91xb35KJJQllB; end sePOIYBEAAbt3DPar8jd5F = ({JuEdAzP84rg2g9z7jUH4CD[16], JuEdAzP84rg2g9z7jUH4CD[16:1]}) + $signed({1'b0, JuEdAzP84rg2g9z7jUH4CD[0]}); iR0ShkyVRkHalUKTDnP0tG = sePOIYBEAAbt3DPar8jd5F >>> 8'd1; j3ureEigNPclVAPr6VwHVbG = {iR0ShkyVRkHalUKTDnP0tG[15:0], 1'b0}; A5SQIaNgqW7DcTqQkKRVeD = j3ureEigNPclVAPr6VwHVbG[15:0]; PmhJP7JCYGM2OStQXGIHgD = ({w13lDdnHeKbz12RPLclXaYB[16], w13lDdnHeKbz12RPLclXaYB[16:1]}) + $signed({1'b0, w13lDdnHeKbz12RPLclXaYB[0]}); TqfF3Zgxtm2cKWvwqij3m = PmhJP7JCYGM2OStQXGIHgD >>> 8'd1; xijHKILnnZ8AgezrLRQvfF = {TqfF3Zgxtm2cKWvwqij3m[15:0], 1'b0}; GaetbCaMty7UkzjqNoYErC = xijHKILnnZ8AgezrLRQvfF[15:0]; LoYaOvLnEQPAYlYtjywSTF = ({G1cI3X0rnsuzwQl9n17YG[16], G1cI3X0rnsuzwQl9n17YG[16:1]}) + $signed({1'b0, G1cI3X0rnsuzwQl9n17YG[0]}); Wf2SXd0xW1vBpZ49DhpQPE = LoYaOvLnEQPAYlYtjywSTF >>> 8'd1; q5X9uuOdY7IBIroLr9svCOD = {Wf2SXd0xW1vBpZ49DhpQPE[15:0], 1'b0}; M5AqS9R7rFTkWxwo8io2rH = q5X9uuOdY7IBIroLr9svCOD[15:0]; BWK9w55Ml1WM8fecaddoXH = ({GXg6LN8xFsDjdENYEDgKvC[16], GXg6LN8xFsDjdENYEDgKvC[16:1]}) + $signed({1'b0, GXg6LN8xFsDjdENYEDgKvC[0]}); h5B5oTxicZ5M23LhruZny = BWK9w55Ml1WM8fecaddoXH >>> 8'd1; DZuRxUKTwIbTxoU1h9ItHG = {h5B5oTxicZ5M23LhruZny[15:0], 1'b0}; lcJo4MnEaj41ofRAtLkn4D = DZuRxUKTwIbTxoU1h9ItHG[15:0]; xijMuK2nBHoByB8rlrH50E = c4yitNmVtLmJQVcYGJPLIKF; end assign B58twvtfgVWGK5P29KavtH = A5SQIaNgqW7DcTqQkKRVeD; assign qhk6Uhwhppvpssqm7Nh6XE = GaetbCaMty7UkzjqNoYErC; assign k3VfrgkD6DWITJL9WW5W4D = M5AqS9R7rFTkWxwo8io2rH; assign pPn6MVGqBLqJ0xzN2WYfFG = lcJo4MnEaj41ofRAtLkn4D; assign jNZ4xylBKAANfCL11XNxzB = xijMuK2nBHoByB8rlrH50E; endmodule