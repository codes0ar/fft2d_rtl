`timescale 1 ns / 1 ns module zVydWOLm2SZCpbjeNcZUmC (v04pHKxyc2sPW047bbyUgE, QDJhCuX1glwonJutj0sIMH, g0hVqHZpe6H7t41TOVwtoTE, qmEenX2Yt9VTzGvbielz5B, DiF2KV4VbJn3P66sh0MYvH, ds3UaO1QhyfiWT7RZKX23G, tCCvu1nsVn6k0oKnEbNi9E); parameter integer AddrWidth = 1; parameter integer DataWidth = 1; input v04pHKxyc2sPW047bbyUgE; input signed [DataWidth - 1:0] QDJhCuX1glwonJutj0sIMH; input signed [DataWidth - 1:0] g0hVqHZpe6H7t41TOVwtoTE; input [AddrWidth - 1:0] qmEenX2Yt9VTzGvbielz5B; input DiF2KV4VbJn3P66sh0MYvH; output signed [DataWidth - 1:0] ds3UaO1QhyfiWT7RZKX23G; output signed [DataWidth - 1:0] tCCvu1nsVn6k0oKnEbNi9E; reg [DataWidth*2 - 1:0] ram [2**AddrWidth - 1:0]; reg [DataWidth*2 - 1:0] data_int; wire cYnz1pueoZwFln8h5mrvmC; always @(posedge v04pHKxyc2sPW047bbyUgE) begin : zVydWOLm2SZCpbjeNcZUmC_prc if (DiF2KV4VbJn3P66sh0MYvH == 1'b1) begin ram[qmEenX2Yt9VTzGvbielz5B] <= {QDJhCuX1glwonJutj0sIMH, g0hVqHZpe6H7t41TOVwtoTE}; data_int <= {QDJhCuX1glwonJutj0sIMH, g0hVqHZpe6H7t41TOVwtoTE}; end else begin data_int <= ram[qmEenX2Yt9VTzGvbielz5B]; end end assign ds3UaO1QhyfiWT7RZKX23G = data_int[DataWidth*2-1:DataWidth]; assign tCCvu1nsVn6k0oKnEbNi9E = data_int[DataWidth-1:0]; endmodule