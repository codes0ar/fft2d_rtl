`timescale 1 ns / 1 ns module xbcMJDB8htpX3R9YnKkaXC (QQYO9noW2AzWAhLJIl3WIE, LIf9KkhuVKSu7vlUpWufBG, c9WUZlfywHR3RaGJnbumYHB, iU3uCiDXuU6z4nkTQ5PufE, z8dRITT2PceChhB9z9EWBC, N7ZKCQ4vfkUB2KkHwgE4GC, PfPBxRXyGunZRp8BSw7dcF, o5kjnQ9W5HT05kz0swOA6QH); input [31:0] QQYO9noW2AzWAhLJIl3WIE; input [31:0] LIf9KkhuVKSu7vlUpWufBG; input [31:0] c9WUZlfywHR3RaGJnbumYHB; input [31:0] iU3uCiDXuU6z4nkTQ5PufE; output [15:0] z8dRITT2PceChhB9z9EWBC; output [15:0] N7ZKCQ4vfkUB2KkHwgE4GC; output [15:0] PfPBxRXyGunZRp8BSw7dcF; output [15:0] o5kjnQ9W5HT05kz0swOA6QH; wire [31:0] yQNwAzareGOhTeFAcGgFWE [0:3]; wire [15:0] sBKdfayBUR3Ntuy7EQrBgD [0:3]; wire [15:0] mOhSSytk7nWnNPtZQ4VYl [0:3]; wire [15:0] Qs9FrBdvqkfYe6HDuZ5x4G [0:3]; wire [15:0] KeIx4znJ7NwHTA7mczkoe [0:3]; wire [15:0] pdFb2Ar1wmoFWvU07SJWFF [0:3]; wire [15:0] QPMLNVTOMA3OrhKJ2KbGiH [0:3]; wire [15:0] DFkPjhhRCMOYOsSbu6aQEF [0:3]; wire [15:0] NtHjaHzNt0xelhyuxLFDIE [0:3]; wire [15:0] vYbET88zhkForoawWcw18E [0:3]; wire [15:0] x1hHF4Y8ZceMfdfnAWH8Mc [0:3]; wire [15:0] Euq2kmsb9LTNk8IgXS0ol [0:3]; wire [15:0] s3eHG7L1MH98LfVKO4py88F [0:3]; wire [15:0] JBmdc6zOYDzlxqcx1YjZb [0:3]; wire [15:0] zawXB1WtJmMfC1cNcABaaE [0:3]; wire [15:0] nORSkpKN0CGUenzeTFfUDB [0:3]; wire [0:3] fXtzdo4P9yi1Ciqp6QBfjC; wire [15:0] ajv4lpvFjoE3ofDGMFu5cE [0:3]; wire [15:0] fatWyfdkxQ7BzaNjbRT4QD [0:3]; wire [0:3] n7hoWcccdXrFN0C874HrpEB; wire [1:0] ebKSCnB4aCunFgmKuqoZYH; wire [1:0] YetQ2qzSWwynIKaYyCEtpC; wire [1:0] vF7LrwtznLIhBcugoROF9E; wire [1:0] EQrAbv0nHPKWlNwGxFRE9; wire [15:0] GySsTihj2cPCBENEuIyCSD [0:3]; wire [15:0] xkbuOVpB2WYtI1blvBLI4F [0:3]; wire [0:3] K3vG6BZkHRRw0KY26D9MZB; wire [1:0] lUScGnUZMrmRi9dRMz0LkD; wire [1:0] TIelA9H027HmZsaaQAWkHE; wire [1:0] TvQBVOfXbi9bTFlCx2e1lD; wire [1:0] s9b257LtpWdWk98ZP3IqF2C; wire [15:0] SrrYc2LpbOfxe2q5vcN0ZB [0:3]; wire [15:0] HXKQBF1mrJNaqSvHX0NNjE [0:3]; wire [0:3] n9yUlIfpQp88T4XdCnh7CDF; wire [1:0] d5CXluM5YmRNluM6LdzEuRD; wire [1:0] MWRVmHwNJJTFsuBNccXpwG; wire [1:0] UeFun2KVGdW93kVlfBFPhD; wire [1:0] EnoEIA9Z5jPxqZoHjfSYbC; wire [15:0] NEJXc3NqgfPBnBXZhsnaBH [0:3]; wire [15:0] pfAEfAzOvu7FtEVFulxbzD [0:3]; wire [0:3] JlM61doAjTFQp2IhAs1cSH; wire [1:0] gBkF6hCOJWWy5LuZbB48v; wire [1:0] aVVNtXP6Zhxq1mxzswY6dD; wire [1:0] lXw2p556JisxQQ4a3indQH; wire [1:0] eMgSW0lzEQfeq7vx5kbytC; wire [15:0] Ndwbn1qn70dbIKd1eeGFLH [0:3]; wire [15:0] w5i8Ug2h8McUnQb3WOIwnOC [0:3]; wire [0:3] yyuLRu89eNc5LwJryJc7rE; wire [1:0] gjjq7XRjRpkPoRKYu5l6n; wire [1:0] hvpZkEPsH8kWqLanUTpxMB; wire [1:0] zmbkHL82PolXRAHTmnIS9D; wire [1:0] g9yIixLFTxnivPa0KqVeY1D; wire [15:0] A4JsqN6vYZ3AEKxV7Ife2D [0:3]; wire [15:0] jqLr7Qvd3gtCcUpcnS2jjE [0:3]; wire [0:3] ScrD9UeAxKjITzyoNx94zC; wire [1:0] ATVtgjciSvCRUI7H3Y9tuD; wire [1:0] w5ir8YG7fu0QbjBpBkweN4; wire [1:0] HWg9kb19eJgbRWUdQ19fQH; wire [1:0] xkG7Las3P9GdNkm3ZSDvCH; wire [15:0] kPPlhFE2ldEEQzJYYPeCpC [0:3]; wire [15:0] f1vtztaLG8k7ETvXjGQi2D [0:3]; wire [0:3] WM76Z8aHuuoFAdf9WffSUE; wire [1:0] FBdqgz94a8SGX1FULhpnhF; wire [1:0] MbKdiATHU4k8jUyFDfh7qF; wire [1:0] eIVteNEy2TzDzIZaAntJEE; wire [1:0] DL0fzBiiKkI4abOA2mryHG; wire [15:0] eq6ExCvRAypD8ZXX1hJg2G [0:3]; wire [15:0] zqoHGtfy6Sfo7Yl3f754XE [0:3]; wire [0:3] TkIpU7Kfy1Dc33ZRJQj19C; wire [1:0] NtsaMyVZXVYmztcjOvOk8; wire [1:0] Ow2gCZKYLWzsXB6jHnoqfG; wire [1:0] otv4IxbTPpKKTvscHxftHG; wire [1:0] l0guWc0JIHa1f8SBb77OlIC; wire [15:0] e1s8qm2TAAcsGxoTmde7BD [0:3]; wire [15:0] PhcezgX6tOzisplfkIJwjD [0:3]; wire [0:3] a99cv4QPwIifb55QksH05aG; wire [1:0] q26YIydocFfUg15Xj6RX5F; wire [1:0] E1ItsZZHtdvolvnwfPb6NC; wire [1:0] PnPVhqoxV0gkaQbzZXf7AD; wire [1:0] n9HtzElTizPjcECkLfcWMT; wire [15:0] N3LfeWGStZMqNRoOruJiLB [0:3]; wire [15:0] Rzd2KleDteHJnQGGQBspBG [0:3]; wire [0:3] rvf3v0TbKi0SUQyjoMm0WE; wire [1:0] K2KmCTF5G7ost89y9oqLiD; wire [1:0] AIcGcubjt3yRVo2TP54CyG; wire [1:0] DPfpo6Ze4IPKLEjjyJWtJD; wire [1:0] DKFv0pTB8YURDrEOItHrZH; wire [15:0] c1ronCM2H01cjuP1wRFxc7C [0:3]; wire [15:0] ue4zD618Z3SRCgWU1P9vMG [0:3]; wire [0:3] M9E8thmcmP8jFioTvkEhuB; wire [1:0] iUgDeFg7wK7VmcsUejECJE; wire [1:0] o6J8Fasm5DBKwavuQUf8xIE; wire [1:0] IqP61QTzblzhrmpI3gXwDD; wire [1:0] LBeizRxhVhpzPZf9SPe9jB; wire [15:0] TKuu61vVE7qT0QqU65DVCB [0:3]; wire [15:0] h75JuQ3GzF4Eyf7QEyVL2ND [0:3]; wire [0:3] taujhy7mQH8DNG1xOnzviE; wire [1:0] CzuyViL53TclNSqIDzrvkF; wire [1:0] p4YcTlbohONe137ErNOKTLG; wire [1:0] H0sU7VFpqA2INbTk7cMsZ; wire [1:0] i9pK5LFhFYyxV7eDKr9g3FD; wire [15:0] UXVpiMug8SwGCNbjOrLnFH [0:3]; wire [15:0] AdUKfM0WY49g0VXTwB2VgF [0:3]; wire hlBwt15h00wuxdBNH1KMDG; assign yQNwAzareGOhTeFAcGgFWE[0] = QQYO9noW2AzWAhLJIl3WIE; assign yQNwAzareGOhTeFAcGgFWE[1] = LIf9KkhuVKSu7vlUpWufBG; assign yQNwAzareGOhTeFAcGgFWE[2] = c9WUZlfywHR3RaGJnbumYHB; assign yQNwAzareGOhTeFAcGgFWE[3] = iU3uCiDXuU6z4nkTQ5PufE; assign sBKdfayBUR3Ntuy7EQrBgD[0] = yQNwAzareGOhTeFAcGgFWE[0][15:0]; assign sBKdfayBUR3Ntuy7EQrBgD[1] = yQNwAzareGOhTeFAcGgFWE[1][15:0]; assign sBKdfayBUR3Ntuy7EQrBgD[2] = yQNwAzareGOhTeFAcGgFWE[2][15:0]; assign sBKdfayBUR3Ntuy7EQrBgD[3] = yQNwAzareGOhTeFAcGgFWE[3][15:0]; assign mOhSSytk7nWnNPtZQ4VYl[0] = 16'b0001000000000000; assign mOhSSytk7nWnNPtZQ4VYl[1] = 16'b0001000000000000; assign mOhSSytk7nWnNPtZQ4VYl[2] = 16'b0001000000000000; assign mOhSSytk7nWnNPtZQ4VYl[3] = 16'b0001000000000000; assign Qs9FrBdvqkfYe6HDuZ5x4G[0] = 16'b0000100000000000; assign Qs9FrBdvqkfYe6HDuZ5x4G[1] = 16'b0000100000000000; assign Qs9FrBdvqkfYe6HDuZ5x4G[2] = 16'b0000100000000000; assign Qs9FrBdvqkfYe6HDuZ5x4G[3] = 16'b0000100000000000; assign KeIx4znJ7NwHTA7mczkoe[0] = 16'b0000010000000000; assign KeIx4znJ7NwHTA7mczkoe[1] = 16'b0000010000000000; assign KeIx4znJ7NwHTA7mczkoe[2] = 16'b0000010000000000; assign KeIx4znJ7NwHTA7mczkoe[3] = 16'b0000010000000000; assign pdFb2Ar1wmoFWvU07SJWFF[0] = 16'b0000001000000000; assign pdFb2Ar1wmoFWvU07SJWFF[1] = 16'b0000001000000000; assign pdFb2Ar1wmoFWvU07SJWFF[2] = 16'b0000001000000000; assign pdFb2Ar1wmoFWvU07SJWFF[3] = 16'b0000001000000000; assign QPMLNVTOMA3OrhKJ2KbGiH[0] = 16'b0000000100000000; assign QPMLNVTOMA3OrhKJ2KbGiH[1] = 16'b0000000100000000; assign QPMLNVTOMA3OrhKJ2KbGiH[2] = 16'b0000000100000000; assign QPMLNVTOMA3OrhKJ2KbGiH[3] = 16'b0000000100000000; assign DFkPjhhRCMOYOsSbu6aQEF[0] = 16'b0000000010000000; assign DFkPjhhRCMOYOsSbu6aQEF[1] = 16'b0000000010000000; assign DFkPjhhRCMOYOsSbu6aQEF[2] = 16'b0000000010000000; assign DFkPjhhRCMOYOsSbu6aQEF[3] = 16'b0000000010000000; assign NtHjaHzNt0xelhyuxLFDIE[0] = 16'b0000000001000000; assign NtHjaHzNt0xelhyuxLFDIE[1] = 16'b0000000001000000; assign NtHjaHzNt0xelhyuxLFDIE[2] = 16'b0000000001000000; assign NtHjaHzNt0xelhyuxLFDIE[3] = 16'b0000000001000000; assign vYbET88zhkForoawWcw18E[0] = 16'b0000000000100000; assign vYbET88zhkForoawWcw18E[1] = 16'b0000000000100000; assign vYbET88zhkForoawWcw18E[2] = 16'b0000000000100000; assign vYbET88zhkForoawWcw18E[3] = 16'b0000000000100000; assign x1hHF4Y8ZceMfdfnAWH8Mc[0] = 16'b0000000000010000; assign x1hHF4Y8ZceMfdfnAWH8Mc[1] = 16'b0000000000010000; assign x1hHF4Y8ZceMfdfnAWH8Mc[2] = 16'b0000000000010000; assign x1hHF4Y8ZceMfdfnAWH8Mc[3] = 16'b0000000000010000; assign Euq2kmsb9LTNk8IgXS0ol[0] = 16'b0000000000001000; assign Euq2kmsb9LTNk8IgXS0ol[1] = 16'b0000000000001000; assign Euq2kmsb9LTNk8IgXS0ol[2] = 16'b0000000000001000; assign Euq2kmsb9LTNk8IgXS0ol[3] = 16'b0000000000001000; assign s3eHG7L1MH98LfVKO4py88F[0] = 16'b0000000000000100; assign s3eHG7L1MH98LfVKO4py88F[1] = 16'b0000000000000100; assign s3eHG7L1MH98LfVKO4py88F[2] = 16'b0000000000000100; assign s3eHG7L1MH98LfVKO4py88F[3] = 16'b0000000000000100; assign JBmdc6zOYDzlxqcx1YjZb[0] = 16'b0000000000000010; assign JBmdc6zOYDzlxqcx1YjZb[1] = 16'b0000000000000010; assign JBmdc6zOYDzlxqcx1YjZb[2] = 16'b0000000000000010; assign JBmdc6zOYDzlxqcx1YjZb[3] = 16'b0000000000000010; assign zawXB1WtJmMfC1cNcABaaE[0] = 16'b0000000000000001; assign zawXB1WtJmMfC1cNcABaaE[1] = 16'b0000000000000001; assign zawXB1WtJmMfC1cNcABaaE[2] = 16'b0000000000000001; assign zawXB1WtJmMfC1cNcABaaE[3] = 16'b0000000000000001; assign nORSkpKN0CGUenzeTFfUDB[0] = sBKdfayBUR3Ntuy7EQrBgD[0] & mOhSSytk7nWnNPtZQ4VYl[0]; assign nORSkpKN0CGUenzeTFfUDB[1] = sBKdfayBUR3Ntuy7EQrBgD[1] & mOhSSytk7nWnNPtZQ4VYl[1]; assign nORSkpKN0CGUenzeTFfUDB[2] = sBKdfayBUR3Ntuy7EQrBgD[2] & mOhSSytk7nWnNPtZQ4VYl[2]; assign nORSkpKN0CGUenzeTFfUDB[3] = sBKdfayBUR3Ntuy7EQrBgD[3] & mOhSSytk7nWnNPtZQ4VYl[3]; assign fXtzdo4P9yi1Ciqp6QBfjC[0] = (|nORSkpKN0CGUenzeTFfUDB[0][15:0]); assign fXtzdo4P9yi1Ciqp6QBfjC[1] = (|nORSkpKN0CGUenzeTFfUDB[1][15:0]); assign fXtzdo4P9yi1Ciqp6QBfjC[2] = (|nORSkpKN0CGUenzeTFfUDB[2][15:0]); assign fXtzdo4P9yi1Ciqp6QBfjC[3] = (|nORSkpKN0CGUenzeTFfUDB[3][15:0]); assign ajv4lpvFjoE3ofDGMFu5cE[0] = {15'b0, fXtzdo4P9yi1Ciqp6QBfjC[0]}; assign ajv4lpvFjoE3ofDGMFu5cE[1] = {15'b0, fXtzdo4P9yi1Ciqp6QBfjC[1]}; assign ajv4lpvFjoE3ofDGMFu5cE[2] = {15'b0, fXtzdo4P9yi1Ciqp6QBfjC[2]}; assign ajv4lpvFjoE3ofDGMFu5cE[3] = {15'b0, fXtzdo4P9yi1Ciqp6QBfjC[3]}; assign fatWyfdkxQ7BzaNjbRT4QD[0] = sBKdfayBUR3Ntuy7EQrBgD[0] & Qs9FrBdvqkfYe6HDuZ5x4G[0]; assign fatWyfdkxQ7BzaNjbRT4QD[1] = sBKdfayBUR3Ntuy7EQrBgD[1] & Qs9FrBdvqkfYe6HDuZ5x4G[1]; assign fatWyfdkxQ7BzaNjbRT4QD[2] = sBKdfayBUR3Ntuy7EQrBgD[2] & Qs9FrBdvqkfYe6HDuZ5x4G[2]; assign fatWyfdkxQ7BzaNjbRT4QD[3] = sBKdfayBUR3Ntuy7EQrBgD[3] & Qs9FrBdvqkfYe6HDuZ5x4G[3]; assign n7hoWcccdXrFN0C874HrpEB[0] = (|fatWyfdkxQ7BzaNjbRT4QD[0][15:0]); assign n7hoWcccdXrFN0C874HrpEB[1] = (|fatWyfdkxQ7BzaNjbRT4QD[1][15:0]); assign n7hoWcccdXrFN0C874HrpEB[2] = (|fatWyfdkxQ7BzaNjbRT4QD[2][15:0]); assign n7hoWcccdXrFN0C874HrpEB[3] = (|fatWyfdkxQ7BzaNjbRT4QD[3][15:0]); assign ebKSCnB4aCunFgmKuqoZYH = {1'b0, n7hoWcccdXrFN0C874HrpEB[0]}; assign GySsTihj2cPCBENEuIyCSD[0] = {13'b0, {ebKSCnB4aCunFgmKuqoZYH, 1'b0}}; assign YetQ2qzSWwynIKaYyCEtpC = {1'b0, n7hoWcccdXrFN0C874HrpEB[1]}; assign GySsTihj2cPCBENEuIyCSD[1] = {13'b0, {YetQ2qzSWwynIKaYyCEtpC, 1'b0}}; assign vF7LrwtznLIhBcugoROF9E = {1'b0, n7hoWcccdXrFN0C874HrpEB[2]}; assign GySsTihj2cPCBENEuIyCSD[2] = {13'b0, {vF7LrwtznLIhBcugoROF9E, 1'b0}}; assign EQrAbv0nHPKWlNwGxFRE9 = {1'b0, n7hoWcccdXrFN0C874HrpEB[3]}; assign GySsTihj2cPCBENEuIyCSD[3] = {13'b0, {EQrAbv0nHPKWlNwGxFRE9, 1'b0}}; assign xkbuOVpB2WYtI1blvBLI4F[0] = sBKdfayBUR3Ntuy7EQrBgD[0] & KeIx4znJ7NwHTA7mczkoe[0]; assign xkbuOVpB2WYtI1blvBLI4F[1] = sBKdfayBUR3Ntuy7EQrBgD[1] & KeIx4znJ7NwHTA7mczkoe[1]; assign xkbuOVpB2WYtI1blvBLI4F[2] = sBKdfayBUR3Ntuy7EQrBgD[2] & KeIx4znJ7NwHTA7mczkoe[2]; assign xkbuOVpB2WYtI1blvBLI4F[3] = sBKdfayBUR3Ntuy7EQrBgD[3] & KeIx4znJ7NwHTA7mczkoe[3]; assign K3vG6BZkHRRw0KY26D9MZB[0] = (|xkbuOVpB2WYtI1blvBLI4F[0][15:0]); assign K3vG6BZkHRRw0KY26D9MZB[1] = (|xkbuOVpB2WYtI1blvBLI4F[1][15:0]); assign K3vG6BZkHRRw0KY26D9MZB[2] = (|xkbuOVpB2WYtI1blvBLI4F[2][15:0]); assign K3vG6BZkHRRw0KY26D9MZB[3] = (|xkbuOVpB2WYtI1blvBLI4F[3][15:0]); assign lUScGnUZMrmRi9dRMz0LkD = {1'b0, K3vG6BZkHRRw0KY26D9MZB[0]}; assign SrrYc2LpbOfxe2q5vcN0ZB[0] = {12'b0, {lUScGnUZMrmRi9dRMz0LkD, 2'b00}}; assign TIelA9H027HmZsaaQAWkHE = {1'b0, K3vG6BZkHRRw0KY26D9MZB[1]}; assign SrrYc2LpbOfxe2q5vcN0ZB[1] = {12'b0, {TIelA9H027HmZsaaQAWkHE, 2'b00}}; assign TvQBVOfXbi9bTFlCx2e1lD = {1'b0, K3vG6BZkHRRw0KY26D9MZB[2]}; assign SrrYc2LpbOfxe2q5vcN0ZB[2] = {12'b0, {TvQBVOfXbi9bTFlCx2e1lD, 2'b00}}; assign s9b257LtpWdWk98ZP3IqF2C = {1'b0, K3vG6BZkHRRw0KY26D9MZB[3]}; assign SrrYc2LpbOfxe2q5vcN0ZB[3] = {12'b0, {s9b257LtpWdWk98ZP3IqF2C, 2'b00}}; assign HXKQBF1mrJNaqSvHX0NNjE[0] = sBKdfayBUR3Ntuy7EQrBgD[0] & pdFb2Ar1wmoFWvU07SJWFF[0]; assign HXKQBF1mrJNaqSvHX0NNjE[1] = sBKdfayBUR3Ntuy7EQrBgD[1] & pdFb2Ar1wmoFWvU07SJWFF[1]; assign HXKQBF1mrJNaqSvHX0NNjE[2] = sBKdfayBUR3Ntuy7EQrBgD[2] & pdFb2Ar1wmoFWvU07SJWFF[2]; assign HXKQBF1mrJNaqSvHX0NNjE[3] = sBKdfayBUR3Ntuy7EQrBgD[3] & pdFb2Ar1wmoFWvU07SJWFF[3]; assign n9yUlIfpQp88T4XdCnh7CDF[0] = (|HXKQBF1mrJNaqSvHX0NNjE[0][15:0]); assign n9yUlIfpQp88T4XdCnh7CDF[1] = (|HXKQBF1mrJNaqSvHX0NNjE[1][15:0]); assign n9yUlIfpQp88T4XdCnh7CDF[2] = (|HXKQBF1mrJNaqSvHX0NNjE[2][15:0]); assign n9yUlIfpQp88T4XdCnh7CDF[3] = (|HXKQBF1mrJNaqSvHX0NNjE[3][15:0]); assign d5CXluM5YmRNluM6LdzEuRD = {1'b0, n9yUlIfpQp88T4XdCnh7CDF[0]}; assign NEJXc3NqgfPBnBXZhsnaBH[0] = {11'b0, {d5CXluM5YmRNluM6LdzEuRD, 3'b000}}; assign MWRVmHwNJJTFsuBNccXpwG = {1'b0, n9yUlIfpQp88T4XdCnh7CDF[1]}; assign NEJXc3NqgfPBnBXZhsnaBH[1] = {11'b0, {MWRVmHwNJJTFsuBNccXpwG, 3'b000}}; assign UeFun2KVGdW93kVlfBFPhD = {1'b0, n9yUlIfpQp88T4XdCnh7CDF[2]}; assign NEJXc3NqgfPBnBXZhsnaBH[2] = {11'b0, {UeFun2KVGdW93kVlfBFPhD, 3'b000}}; assign EnoEIA9Z5jPxqZoHjfSYbC = {1'b0, n9yUlIfpQp88T4XdCnh7CDF[3]}; assign NEJXc3NqgfPBnBXZhsnaBH[3] = {11'b0, {EnoEIA9Z5jPxqZoHjfSYbC, 3'b000}}; assign pfAEfAzOvu7FtEVFulxbzD[0] = sBKdfayBUR3Ntuy7EQrBgD[0] & QPMLNVTOMA3OrhKJ2KbGiH[0]; assign pfAEfAzOvu7FtEVFulxbzD[1] = sBKdfayBUR3Ntuy7EQrBgD[1] & QPMLNVTOMA3OrhKJ2KbGiH[1]; assign pfAEfAzOvu7FtEVFulxbzD[2] = sBKdfayBUR3Ntuy7EQrBgD[2] & QPMLNVTOMA3OrhKJ2KbGiH[2]; assign pfAEfAzOvu7FtEVFulxbzD[3] = sBKdfayBUR3Ntuy7EQrBgD[3] & QPMLNVTOMA3OrhKJ2KbGiH[3]; assign JlM61doAjTFQp2IhAs1cSH[0] = (|pfAEfAzOvu7FtEVFulxbzD[0][15:0]); assign JlM61doAjTFQp2IhAs1cSH[1] = (|pfAEfAzOvu7FtEVFulxbzD[1][15:0]); assign JlM61doAjTFQp2IhAs1cSH[2] = (|pfAEfAzOvu7FtEVFulxbzD[2][15:0]); assign JlM61doAjTFQp2IhAs1cSH[3] = (|pfAEfAzOvu7FtEVFulxbzD[3][15:0]); assign gBkF6hCOJWWy5LuZbB48v = {1'b0, JlM61doAjTFQp2IhAs1cSH[0]}; assign Ndwbn1qn70dbIKd1eeGFLH[0] = {10'b0, {gBkF6hCOJWWy5LuZbB48v, 4'b0000}}; assign aVVNtXP6Zhxq1mxzswY6dD = {1'b0, JlM61doAjTFQp2IhAs1cSH[1]}; assign Ndwbn1qn70dbIKd1eeGFLH[1] = {10'b0, {aVVNtXP6Zhxq1mxzswY6dD, 4'b0000}}; assign lXw2p556JisxQQ4a3indQH = {1'b0, JlM61doAjTFQp2IhAs1cSH[2]}; assign Ndwbn1qn70dbIKd1eeGFLH[2] = {10'b0, {lXw2p556JisxQQ4a3indQH, 4'b0000}}; assign eMgSW0lzEQfeq7vx5kbytC = {1'b0, JlM61doAjTFQp2IhAs1cSH[3]}; assign Ndwbn1qn70dbIKd1eeGFLH[3] = {10'b0, {eMgSW0lzEQfeq7vx5kbytC, 4'b0000}}; assign w5i8Ug2h8McUnQb3WOIwnOC[0] = sBKdfayBUR3Ntuy7EQrBgD[0] & DFkPjhhRCMOYOsSbu6aQEF[0]; assign w5i8Ug2h8McUnQb3WOIwnOC[1] = sBKdfayBUR3Ntuy7EQrBgD[1] & DFkPjhhRCMOYOsSbu6aQEF[1]; assign w5i8Ug2h8McUnQb3WOIwnOC[2] = sBKdfayBUR3Ntuy7EQrBgD[2] & DFkPjhhRCMOYOsSbu6aQEF[2]; assign w5i8Ug2h8McUnQb3WOIwnOC[3] = sBKdfayBUR3Ntuy7EQrBgD[3] & DFkPjhhRCMOYOsSbu6aQEF[3]; assign yyuLRu89eNc5LwJryJc7rE[0] = (|w5i8Ug2h8McUnQb3WOIwnOC[0][15:0]); assign yyuLRu89eNc5LwJryJc7rE[1] = (|w5i8Ug2h8McUnQb3WOIwnOC[1][15:0]); assign yyuLRu89eNc5LwJryJc7rE[2] = (|w5i8Ug2h8McUnQb3WOIwnOC[2][15:0]); assign yyuLRu89eNc5LwJryJc7rE[3] = (|w5i8Ug2h8McUnQb3WOIwnOC[3][15:0]); assign gjjq7XRjRpkPoRKYu5l6n = {1'b0, yyuLRu89eNc5LwJryJc7rE[0]}; assign A4JsqN6vYZ3AEKxV7Ife2D[0] = {9'b0, {gjjq7XRjRpkPoRKYu5l6n, 5'b00000}}; assign hvpZkEPsH8kWqLanUTpxMB = {1'b0, yyuLRu89eNc5LwJryJc7rE[1]}; assign A4JsqN6vYZ3AEKxV7Ife2D[1] = {9'b0, {hvpZkEPsH8kWqLanUTpxMB, 5'b00000}}; assign zmbkHL82PolXRAHTmnIS9D = {1'b0, yyuLRu89eNc5LwJryJc7rE[2]}; assign A4JsqN6vYZ3AEKxV7Ife2D[2] = {9'b0, {zmbkHL82PolXRAHTmnIS9D, 5'b00000}}; assign g9yIixLFTxnivPa0KqVeY1D = {1'b0, yyuLRu89eNc5LwJryJc7rE[3]}; assign A4JsqN6vYZ3AEKxV7Ife2D[3] = {9'b0, {g9yIixLFTxnivPa0KqVeY1D, 5'b00000}}; assign jqLr7Qvd3gtCcUpcnS2jjE[0] = sBKdfayBUR3Ntuy7EQrBgD[0] & NtHjaHzNt0xelhyuxLFDIE[0]; assign jqLr7Qvd3gtCcUpcnS2jjE[1] = sBKdfayBUR3Ntuy7EQrBgD[1] & NtHjaHzNt0xelhyuxLFDIE[1]; assign jqLr7Qvd3gtCcUpcnS2jjE[2] = sBKdfayBUR3Ntuy7EQrBgD[2] & NtHjaHzNt0xelhyuxLFDIE[2]; assign jqLr7Qvd3gtCcUpcnS2jjE[3] = sBKdfayBUR3Ntuy7EQrBgD[3] & NtHjaHzNt0xelhyuxLFDIE[3]; assign ScrD9UeAxKjITzyoNx94zC[0] = (|jqLr7Qvd3gtCcUpcnS2jjE[0][15:0]); assign ScrD9UeAxKjITzyoNx94zC[1] = (|jqLr7Qvd3gtCcUpcnS2jjE[1][15:0]); assign ScrD9UeAxKjITzyoNx94zC[2] = (|jqLr7Qvd3gtCcUpcnS2jjE[2][15:0]); assign ScrD9UeAxKjITzyoNx94zC[3] = (|jqLr7Qvd3gtCcUpcnS2jjE[3][15:0]); assign ATVtgjciSvCRUI7H3Y9tuD = {1'b0, ScrD9UeAxKjITzyoNx94zC[0]}; assign kPPlhFE2ldEEQzJYYPeCpC[0] = {8'b0, {ATVtgjciSvCRUI7H3Y9tuD, 6'b000000}}; assign w5ir8YG7fu0QbjBpBkweN4 = {1'b0, ScrD9UeAxKjITzyoNx94zC[1]}; assign kPPlhFE2ldEEQzJYYPeCpC[1] = {8'b0, {w5ir8YG7fu0QbjBpBkweN4, 6'b000000}}; assign HWg9kb19eJgbRWUdQ19fQH = {1'b0, ScrD9UeAxKjITzyoNx94zC[2]}; assign kPPlhFE2ldEEQzJYYPeCpC[2] = {8'b0, {HWg9kb19eJgbRWUdQ19fQH, 6'b000000}}; assign xkG7Las3P9GdNkm3ZSDvCH = {1'b0, ScrD9UeAxKjITzyoNx94zC[3]}; assign kPPlhFE2ldEEQzJYYPeCpC[3] = {8'b0, {xkG7Las3P9GdNkm3ZSDvCH, 6'b000000}}; assign f1vtztaLG8k7ETvXjGQi2D[0] = sBKdfayBUR3Ntuy7EQrBgD[0] & vYbET88zhkForoawWcw18E[0]; assign f1vtztaLG8k7ETvXjGQi2D[1] = sBKdfayBUR3Ntuy7EQrBgD[1] & vYbET88zhkForoawWcw18E[1]; assign f1vtztaLG8k7ETvXjGQi2D[2] = sBKdfayBUR3Ntuy7EQrBgD[2] & vYbET88zhkForoawWcw18E[2]; assign f1vtztaLG8k7ETvXjGQi2D[3] = sBKdfayBUR3Ntuy7EQrBgD[3] & vYbET88zhkForoawWcw18E[3]; assign WM76Z8aHuuoFAdf9WffSUE[0] = (|f1vtztaLG8k7ETvXjGQi2D[0][15:0]); assign WM76Z8aHuuoFAdf9WffSUE[1] = (|f1vtztaLG8k7ETvXjGQi2D[1][15:0]); assign WM76Z8aHuuoFAdf9WffSUE[2] = (|f1vtztaLG8k7ETvXjGQi2D[2][15:0]); assign WM76Z8aHuuoFAdf9WffSUE[3] = (|f1vtztaLG8k7ETvXjGQi2D[3][15:0]); assign FBdqgz94a8SGX1FULhpnhF = {1'b0, WM76Z8aHuuoFAdf9WffSUE[0]}; assign eq6ExCvRAypD8ZXX1hJg2G[0] = {7'b0, {FBdqgz94a8SGX1FULhpnhF, 7'b0000000}}; assign MbKdiATHU4k8jUyFDfh7qF = {1'b0, WM76Z8aHuuoFAdf9WffSUE[1]}; assign eq6ExCvRAypD8ZXX1hJg2G[1] = {7'b0, {MbKdiATHU4k8jUyFDfh7qF, 7'b0000000}}; assign eIVteNEy2TzDzIZaAntJEE = {1'b0, WM76Z8aHuuoFAdf9WffSUE[2]}; assign eq6ExCvRAypD8ZXX1hJg2G[2] = {7'b0, {eIVteNEy2TzDzIZaAntJEE, 7'b0000000}}; assign DL0fzBiiKkI4abOA2mryHG = {1'b0, WM76Z8aHuuoFAdf9WffSUE[3]}; assign eq6ExCvRAypD8ZXX1hJg2G[3] = {7'b0, {DL0fzBiiKkI4abOA2mryHG, 7'b0000000}}; assign zqoHGtfy6Sfo7Yl3f754XE[0] = sBKdfayBUR3Ntuy7EQrBgD[0] & x1hHF4Y8ZceMfdfnAWH8Mc[0]; assign zqoHGtfy6Sfo7Yl3f754XE[1] = sBKdfayBUR3Ntuy7EQrBgD[1] & x1hHF4Y8ZceMfdfnAWH8Mc[1]; assign zqoHGtfy6Sfo7Yl3f754XE[2] = sBKdfayBUR3Ntuy7EQrBgD[2] & x1hHF4Y8ZceMfdfnAWH8Mc[2]; assign zqoHGtfy6Sfo7Yl3f754XE[3] = sBKdfayBUR3Ntuy7EQrBgD[3] & x1hHF4Y8ZceMfdfnAWH8Mc[3]; assign TkIpU7Kfy1Dc33ZRJQj19C[0] = (|zqoHGtfy6Sfo7Yl3f754XE[0][15:0]); assign TkIpU7Kfy1Dc33ZRJQj19C[1] = (|zqoHGtfy6Sfo7Yl3f754XE[1][15:0]); assign TkIpU7Kfy1Dc33ZRJQj19C[2] = (|zqoHGtfy6Sfo7Yl3f754XE[2][15:0]); assign TkIpU7Kfy1Dc33ZRJQj19C[3] = (|zqoHGtfy6Sfo7Yl3f754XE[3][15:0]); assign NtsaMyVZXVYmztcjOvOk8 = {1'b0, TkIpU7Kfy1Dc33ZRJQj19C[0]}; assign e1s8qm2TAAcsGxoTmde7BD[0] = {6'b0, {NtsaMyVZXVYmztcjOvOk8, 8'b00000000}}; assign Ow2gCZKYLWzsXB6jHnoqfG = {1'b0, TkIpU7Kfy1Dc33ZRJQj19C[1]}; assign e1s8qm2TAAcsGxoTmde7BD[1] = {6'b0, {Ow2gCZKYLWzsXB6jHnoqfG, 8'b00000000}}; assign otv4IxbTPpKKTvscHxftHG = {1'b0, TkIpU7Kfy1Dc33ZRJQj19C[2]}; assign e1s8qm2TAAcsGxoTmde7BD[2] = {6'b0, {otv4IxbTPpKKTvscHxftHG, 8'b00000000}}; assign l0guWc0JIHa1f8SBb77OlIC = {1'b0, TkIpU7Kfy1Dc33ZRJQj19C[3]}; assign e1s8qm2TAAcsGxoTmde7BD[3] = {6'b0, {l0guWc0JIHa1f8SBb77OlIC, 8'b00000000}}; assign PhcezgX6tOzisplfkIJwjD[0] = sBKdfayBUR3Ntuy7EQrBgD[0] & Euq2kmsb9LTNk8IgXS0ol[0]; assign PhcezgX6tOzisplfkIJwjD[1] = sBKdfayBUR3Ntuy7EQrBgD[1] & Euq2kmsb9LTNk8IgXS0ol[1]; assign PhcezgX6tOzisplfkIJwjD[2] = sBKdfayBUR3Ntuy7EQrBgD[2] & Euq2kmsb9LTNk8IgXS0ol[2]; assign PhcezgX6tOzisplfkIJwjD[3] = sBKdfayBUR3Ntuy7EQrBgD[3] & Euq2kmsb9LTNk8IgXS0ol[3]; assign a99cv4QPwIifb55QksH05aG[0] = (|PhcezgX6tOzisplfkIJwjD[0][15:0]); assign a99cv4QPwIifb55QksH05aG[1] = (|PhcezgX6tOzisplfkIJwjD[1][15:0]); assign a99cv4QPwIifb55QksH05aG[2] = (|PhcezgX6tOzisplfkIJwjD[2][15:0]); assign a99cv4QPwIifb55QksH05aG[3] = (|PhcezgX6tOzisplfkIJwjD[3][15:0]); assign q26YIydocFfUg15Xj6RX5F = {1'b0, a99cv4QPwIifb55QksH05aG[0]}; assign N3LfeWGStZMqNRoOruJiLB[0] = {5'b0, {q26YIydocFfUg15Xj6RX5F, 9'b000000000}}; assign E1ItsZZHtdvolvnwfPb6NC = {1'b0, a99cv4QPwIifb55QksH05aG[1]}; assign N3LfeWGStZMqNRoOruJiLB[1] = {5'b0, {E1ItsZZHtdvolvnwfPb6NC, 9'b000000000}}; assign PnPVhqoxV0gkaQbzZXf7AD = {1'b0, a99cv4QPwIifb55QksH05aG[2]}; assign N3LfeWGStZMqNRoOruJiLB[2] = {5'b0, {PnPVhqoxV0gkaQbzZXf7AD, 9'b000000000}}; assign n9HtzElTizPjcECkLfcWMT = {1'b0, a99cv4QPwIifb55QksH05aG[3]}; assign N3LfeWGStZMqNRoOruJiLB[3] = {5'b0, {n9HtzElTizPjcECkLfcWMT, 9'b000000000}}; assign Rzd2KleDteHJnQGGQBspBG[0] = sBKdfayBUR3Ntuy7EQrBgD[0] & s3eHG7L1MH98LfVKO4py88F[0]; assign Rzd2KleDteHJnQGGQBspBG[1] = sBKdfayBUR3Ntuy7EQrBgD[1] & s3eHG7L1MH98LfVKO4py88F[1]; assign Rzd2KleDteHJnQGGQBspBG[2] = sBKdfayBUR3Ntuy7EQrBgD[2] & s3eHG7L1MH98LfVKO4py88F[2]; assign Rzd2KleDteHJnQGGQBspBG[3] = sBKdfayBUR3Ntuy7EQrBgD[3] & s3eHG7L1MH98LfVKO4py88F[3]; assign rvf3v0TbKi0SUQyjoMm0WE[0] = (|Rzd2KleDteHJnQGGQBspBG[0][15:0]); assign rvf3v0TbKi0SUQyjoMm0WE[1] = (|Rzd2KleDteHJnQGGQBspBG[1][15:0]); assign rvf3v0TbKi0SUQyjoMm0WE[2] = (|Rzd2KleDteHJnQGGQBspBG[2][15:0]); assign rvf3v0TbKi0SUQyjoMm0WE[3] = (|Rzd2KleDteHJnQGGQBspBG[3][15:0]); assign K2KmCTF5G7ost89y9oqLiD = {1'b0, rvf3v0TbKi0SUQyjoMm0WE[0]}; assign c1ronCM2H01cjuP1wRFxc7C[0] = {4'b0, {K2KmCTF5G7ost89y9oqLiD, 10'b0000000000}}; assign AIcGcubjt3yRVo2TP54CyG = {1'b0, rvf3v0TbKi0SUQyjoMm0WE[1]}; assign c1ronCM2H01cjuP1wRFxc7C[1] = {4'b0, {AIcGcubjt3yRVo2TP54CyG, 10'b0000000000}}; assign DPfpo6Ze4IPKLEjjyJWtJD = {1'b0, rvf3v0TbKi0SUQyjoMm0WE[2]}; assign c1ronCM2H01cjuP1wRFxc7C[2] = {4'b0, {DPfpo6Ze4IPKLEjjyJWtJD, 10'b0000000000}}; assign DKFv0pTB8YURDrEOItHrZH = {1'b0, rvf3v0TbKi0SUQyjoMm0WE[3]}; assign c1ronCM2H01cjuP1wRFxc7C[3] = {4'b0, {DKFv0pTB8YURDrEOItHrZH, 10'b0000000000}}; assign ue4zD618Z3SRCgWU1P9vMG[0] = sBKdfayBUR3Ntuy7EQrBgD[0] & JBmdc6zOYDzlxqcx1YjZb[0]; assign ue4zD618Z3SRCgWU1P9vMG[1] = sBKdfayBUR3Ntuy7EQrBgD[1] & JBmdc6zOYDzlxqcx1YjZb[1]; assign ue4zD618Z3SRCgWU1P9vMG[2] = sBKdfayBUR3Ntuy7EQrBgD[2] & JBmdc6zOYDzlxqcx1YjZb[2]; assign ue4zD618Z3SRCgWU1P9vMG[3] = sBKdfayBUR3Ntuy7EQrBgD[3] & JBmdc6zOYDzlxqcx1YjZb[3]; assign M9E8thmcmP8jFioTvkEhuB[0] = (|ue4zD618Z3SRCgWU1P9vMG[0][15:0]); assign M9E8thmcmP8jFioTvkEhuB[1] = (|ue4zD618Z3SRCgWU1P9vMG[1][15:0]); assign M9E8thmcmP8jFioTvkEhuB[2] = (|ue4zD618Z3SRCgWU1P9vMG[2][15:0]); assign M9E8thmcmP8jFioTvkEhuB[3] = (|ue4zD618Z3SRCgWU1P9vMG[3][15:0]); assign iUgDeFg7wK7VmcsUejECJE = {1'b0, M9E8thmcmP8jFioTvkEhuB[0]}; assign TKuu61vVE7qT0QqU65DVCB[0] = {3'b0, {iUgDeFg7wK7VmcsUejECJE, 11'b00000000000}}; assign o6J8Fasm5DBKwavuQUf8xIE = {1'b0, M9E8thmcmP8jFioTvkEhuB[1]}; assign TKuu61vVE7qT0QqU65DVCB[1] = {3'b0, {o6J8Fasm5DBKwavuQUf8xIE, 11'b00000000000}}; assign IqP61QTzblzhrmpI3gXwDD = {1'b0, M9E8thmcmP8jFioTvkEhuB[2]}; assign TKuu61vVE7qT0QqU65DVCB[2] = {3'b0, {IqP61QTzblzhrmpI3gXwDD, 11'b00000000000}}; assign LBeizRxhVhpzPZf9SPe9jB = {1'b0, M9E8thmcmP8jFioTvkEhuB[3]}; assign TKuu61vVE7qT0QqU65DVCB[3] = {3'b0, {LBeizRxhVhpzPZf9SPe9jB, 11'b00000000000}}; assign h75JuQ3GzF4Eyf7QEyVL2ND[0] = sBKdfayBUR3Ntuy7EQrBgD[0] & zawXB1WtJmMfC1cNcABaaE[0]; assign h75JuQ3GzF4Eyf7QEyVL2ND[1] = sBKdfayBUR3Ntuy7EQrBgD[1] & zawXB1WtJmMfC1cNcABaaE[1]; assign h75JuQ3GzF4Eyf7QEyVL2ND[2] = sBKdfayBUR3Ntuy7EQrBgD[2] & zawXB1WtJmMfC1cNcABaaE[2]; assign h75JuQ3GzF4Eyf7QEyVL2ND[3] = sBKdfayBUR3Ntuy7EQrBgD[3] & zawXB1WtJmMfC1cNcABaaE[3]; assign taujhy7mQH8DNG1xOnzviE[0] = (|h75JuQ3GzF4Eyf7QEyVL2ND[0][15:0]); assign taujhy7mQH8DNG1xOnzviE[1] = (|h75JuQ3GzF4Eyf7QEyVL2ND[1][15:0]); assign taujhy7mQH8DNG1xOnzviE[2] = (|h75JuQ3GzF4Eyf7QEyVL2ND[2][15:0]); assign taujhy7mQH8DNG1xOnzviE[3] = (|h75JuQ3GzF4Eyf7QEyVL2ND[3][15:0]); assign CzuyViL53TclNSqIDzrvkF = {1'b0, taujhy7mQH8DNG1xOnzviE[0]}; assign UXVpiMug8SwGCNbjOrLnFH[0] = {2'b0, {CzuyViL53TclNSqIDzrvkF, 12'b000000000000}}; assign p4YcTlbohONe137ErNOKTLG = {1'b0, taujhy7mQH8DNG1xOnzviE[1]}; assign UXVpiMug8SwGCNbjOrLnFH[1] = {2'b0, {p4YcTlbohONe137ErNOKTLG, 12'b000000000000}}; assign H0sU7VFpqA2INbTk7cMsZ = {1'b0, taujhy7mQH8DNG1xOnzviE[2]}; assign UXVpiMug8SwGCNbjOrLnFH[2] = {2'b0, {H0sU7VFpqA2INbTk7cMsZ, 12'b000000000000}}; assign i9pK5LFhFYyxV7eDKr9g3FD = {1'b0, taujhy7mQH8DNG1xOnzviE[3]}; assign UXVpiMug8SwGCNbjOrLnFH[3] = {2'b0, {i9pK5LFhFYyxV7eDKr9g3FD, 12'b000000000000}}; assign AdUKfM0WY49g0VXTwB2VgF[0] = UXVpiMug8SwGCNbjOrLnFH[0] | (TKuu61vVE7qT0QqU65DVCB[0] | (c1ronCM2H01cjuP1wRFxc7C[0] | (N3LfeWGStZMqNRoOruJiLB[0] | (e1s8qm2TAAcsGxoTmde7BD[0] | (eq6ExCvRAypD8ZXX1hJg2G[0] | (kPPlhFE2ldEEQzJYYPeCpC[0] | (A4JsqN6vYZ3AEKxV7Ife2D[0] | (Ndwbn1qn70dbIKd1eeGFLH[0] | (NEJXc3NqgfPBnBXZhsnaBH[0] | (SrrYc2LpbOfxe2q5vcN0ZB[0] | (ajv4lpvFjoE3ofDGMFu5cE[0] | GySsTihj2cPCBENEuIyCSD[0]))))))))))); assign AdUKfM0WY49g0VXTwB2VgF[1] = UXVpiMug8SwGCNbjOrLnFH[1] | (TKuu61vVE7qT0QqU65DVCB[1] | (c1ronCM2H01cjuP1wRFxc7C[1] | (N3LfeWGStZMqNRoOruJiLB[1] | (e1s8qm2TAAcsGxoTmde7BD[1] | (eq6ExCvRAypD8ZXX1hJg2G[1] | (kPPlhFE2ldEEQzJYYPeCpC[1] | (A4JsqN6vYZ3AEKxV7Ife2D[1] | (Ndwbn1qn70dbIKd1eeGFLH[1] | (NEJXc3NqgfPBnBXZhsnaBH[1] | (SrrYc2LpbOfxe2q5vcN0ZB[1] | (ajv4lpvFjoE3ofDGMFu5cE[1] | GySsTihj2cPCBENEuIyCSD[1]))))))))))); assign AdUKfM0WY49g0VXTwB2VgF[2] = UXVpiMug8SwGCNbjOrLnFH[2] | (TKuu61vVE7qT0QqU65DVCB[2] | (c1ronCM2H01cjuP1wRFxc7C[2] | (N3LfeWGStZMqNRoOruJiLB[2] | (e1s8qm2TAAcsGxoTmde7BD[2] | (eq6ExCvRAypD8ZXX1hJg2G[2] | (kPPlhFE2ldEEQzJYYPeCpC[2] | (A4JsqN6vYZ3AEKxV7Ife2D[2] | (Ndwbn1qn70dbIKd1eeGFLH[2] | (NEJXc3NqgfPBnBXZhsnaBH[2] | (SrrYc2LpbOfxe2q5vcN0ZB[2] | (ajv4lpvFjoE3ofDGMFu5cE[2] | GySsTihj2cPCBENEuIyCSD[2]))))))))))); assign AdUKfM0WY49g0VXTwB2VgF[3] = UXVpiMug8SwGCNbjOrLnFH[3] | (TKuu61vVE7qT0QqU65DVCB[3] | (c1ronCM2H01cjuP1wRFxc7C[3] | (N3LfeWGStZMqNRoOruJiLB[3] | (e1s8qm2TAAcsGxoTmde7BD[3] | (eq6ExCvRAypD8ZXX1hJg2G[3] | (kPPlhFE2ldEEQzJYYPeCpC[3] | (A4JsqN6vYZ3AEKxV7Ife2D[3] | (Ndwbn1qn70dbIKd1eeGFLH[3] | (NEJXc3NqgfPBnBXZhsnaBH[3] | (SrrYc2LpbOfxe2q5vcN0ZB[3] | (ajv4lpvFjoE3ofDGMFu5cE[3] | GySsTihj2cPCBENEuIyCSD[3]))))))))))); assign z8dRITT2PceChhB9z9EWBC = AdUKfM0WY49g0VXTwB2VgF[0]; assign N7ZKCQ4vfkUB2KkHwgE4GC = AdUKfM0WY49g0VXTwB2VgF[1]; assign PfPBxRXyGunZRp8BSw7dcF = AdUKfM0WY49g0VXTwB2VgF[2]; assign o5kjnQ9W5HT05kz0swOA6QH = AdUKfM0WY49g0VXTwB2VgF[3]; endmodule