`timescale 1 ns / 1 ns module fft2d (mclk, rstb, qdin_0, qdin_1, qdin_2, qdin_3, f1en, srst, f2Vld, f2abs_0, f2abs_1, f2abs_2, f2abs_3); input mclk; input rstb; input signed [15:0] qdin_0; input signed [15:0] qdin_1; input signed [15:0] qdin_2; input signed [15:0] qdin_3; input f1en; input srst; output f2Vld; output [15:0] f2abs_0; output [15:0] f2abs_1; output [15:0] f2abs_2; output [15:0] f2abs_3; wire signed [15:0] RDoofzNe0oXjNKPxTYnsJG; wire signed [15:0] l96ToZvA3JxZRoamoFQ1UB; wire signed [15:0] vuBZeR1bCIQ7eYub4Nym0B; wire signed [15:0] kYezVXe7e7E7TbchXde4QG; wire signed [15:0] BdTGl8ppsd8fNRyihNQvWD; wire signed [15:0] j5vaJTpXoIQ2WMB1cDQvqC; wire signed [15:0] fijzTATvD4NCVDjSoyqDXC; wire signed [15:0] uH5IsuPlvOkkvGQhI40ZZF; wire TciTCDpCygk823aRzOkhCE; reg [21:0] lYL40DZJNrZGA50HVltAXD; wire [43:0] d5CXluM5YmRNluM6LdzEuRD; wire [17:0] jAqDYspp5RSupfEc9vWoJH; wire HHiAQq0eXS4V724AeWtEMD; wire [16:0] PFHmZS0ipZLKqJ39A27L8F; wire [31:0] HtkwvAWd5V10OAKRmUTiLD; wire [31:0] IMy6yN0h9YqHeUl7378ZhB; wire [63:0] FBdqgz94a8SGX1FULhpnhF; wire [9:0] eq6ExCvRAypD8ZXX1hJg2G; wire [31:0] M6DCmjjEAXTHH63S0PcE0E; wire [15:0] ImRl6qg5Qleo28k6kzf5ID; wire [31:0] xWllAgKkXsJdEckAS1JkRE; wire [16:0] txIZVPOqyNjR0XJaNnEWgC; wire [16:0] o8JfccMcxN3IkRA878Wl6qB [0:3]; wire [16:0] iVUCRzTzoib1t9JQL19F1B [0:3]; wire [1:0] q8UubaExFIU37MrHaKCYjEH [0:3]; wire signed [32:0] i3T8rgFVbtYhLp11xyNVaG; wire signed [32:0] xb5OWtSspXT5QIrsjYRNyC; wire signed [32:0] zkeZd8GIm1z3m743ZzXwoF; wire signed [32:0] d3io0lXPWPHhxjlWak3S1G; wire signed [32:0] kmQDARJ5RSC33fkFkFEZvB [0:3]; wire [63:0] h6X6Ift6lj74yXs2DyR91PG; wire [31:0] v0ZPFDd9cyRidUk0uUpeZF; wire [15:0] UGX8fdfHPAfRuWbIXSAJkC; wire [31:0] iUgDeFg7wK7VmcsUejECJE; wire [16:0] kXQPeGN2PPqOhoBeXJau8E; wire [16:0] RgAX8O9DbR6HNMiXsFyzb [0:3]; wire [16:0] Hm89BMHiz5dcKMTSyT6ZgE [0:3]; wire [1:0] TqEdytxeoETbv4LqQENvdE [0:3]; wire signed [32:0] HWvpOqHBtG8nHbtWWOs5ME [0:3]; wire signed [32:0] XFDR6Vjpsj8y8if8sCJpyC [0:3]; reg signed [32:0] ZIXwDtDHOFCY284ItMUkPE [0:3]; reg wmHZAgpaaD0AnBPdMzFAWB; wire [16:0] JM1PWrdw4CsiaxhIFEj0FG [0:3]; wire [33:0] NtsaMyVZXVYmztcjOvOk8; wire [33:0] Ow2gCZKYLWzsXB6jHnoqfG; wire [33:0] otv4IxbTPpKKTvscHxftHG; wire [33:0] l0guWc0JIHa1f8SBb77OlIC; wire [16:0] Bx5GbZBMMZWJmhJNe1plNE [0:3]; wire [17:0] vDf5jyCbwqHvGEEIH52rqG [0:3]; wire [31:0] KyXrE6JYq7NUB9MlwmKcGH; wire [31:0] THQEaifSmIkcouXcNP6X2G; wire [31:0] Xp7jYGB4wGPVX0g6nIaYOD; wire [15:0] x2T5MHXEjHB4mbeunlQ5xlC; wire [15:0] m3srRE1KQDnmVOjclDlFnB; wire [15:0] cZMBbP0tbfriJB96bWdXBG; wire [15:0] OlmksAU0OqEmB1eHPlD4LF; wire [15:0] wZQ5Nh8v8jyFGZaqm7MPFF [0:3]; wire [31:0] K2KmCTF5G7ost89y9oqLiD; wire [31:0] AIcGcubjt3yRVo2TP54CyG; wire [31:0] DPfpo6Ze4IPKLEjjyJWtJD; wire [31:0] DKFv0pTB8YURDrEOItHrZH; wire [16:0] n7lC0EX54a5Db2Ey78BZWH [0:3]; wire [33:0] gjjq7XRjRpkPoRKYu5l6n; wire [33:0] hvpZkEPsH8kWqLanUTpxMB; wire [33:0] zmbkHL82PolXRAHTmnIS9D; wire [33:0] g9yIixLFTxnivPa0KqVeY1D; wire [16:0] mhinOy8fRr1hyDeV9qCPFB [0:3]; wire [33:0] ATVtgjciSvCRUI7H3Y9tuD; wire [9:0] toucxMaGXtuei4mJhB7SvH; wire [17:0] t1mfqjXjUa0cnuylRz3bBNF; wire [17:0] BQWUnHpxPEGrMvfoEg50BE [0:3]; wire [17:0] UIikZeafI7JRbAIwWZXxZG; wire [17:0] YHsZm9RxIvVHFFCFqjHJbB; wire [17:0] Ro8Qq6Y03XDjqsnyirVcTD; wire [17:0] XW2XizJGnQkUYhMVZ7vzD; wire [17:0] KRGfxNqFr6P3qLzrH4DIYD [0:3]; wire [17:0] YkB06NLyXnKPFxzf13DnpH [0:3]; wire [16:0] gAw9zJNNZqPQfnlAoc3jXH [0:3]; wire signed [15:0] CqX3zbRXkD0JZjUDCE4uyC [0:3]; wire signed [15:0] Y2qRC0lD6WkLUd7tO2DL8D [0:3]; wire signed [15:0] w27urwsxsx3vX1J4eEaqy0D; wire signed [15:0] onEIj0VH5ehJOImYn9CHFC; wire signed [15:0] GyXnWgCHVjevCAC5dsEk8G; wire signed [15:0] dCpVrDZOfokUK9iu0jbwzC; wire signed [15:0] h8Njhoqboql6ktvl74YNlD; wire signed [15:0] g0CmNQp5HtaKwsfnggkLOD; wire signed [15:0] r7YnXgwRbNGWdEl2TZcAw0C; wire signed [15:0] u1xFlD3D83sqzZNknRicP6B; wire signed [15:0] M5pFttxc4QndsuSd89rKrD; wire signed [15:0] FVvSvaFiVsOXZzGo86bsoC; wire signed [15:0] dte5acyHW51RNSwjPM8XJD; wire signed [15:0] wLogEYXttTcYn1hYyKkIwE; wire signed [15:0] Z1XJpcLo4zUnViPcNLmlmC; wire signed [15:0] yfb14sul5mbLBMqiwceCCC; wire signed [15:0] nz8qYIrRTZKfZJZAE7BZrF; wire signed [15:0] iZEHwpNoTE4xYjGNgFVDSH; wire signed [15:0] AvHKfOLcDBK6tGfufEsPhF [0:3]; wire signed [15:0] AUkBI5w4Pfinl5l6Ts0oXB [0:3]; wire [17:0] perQtgyUzTQmgJPDhQgq5D [0:3]; wire [17:0] wnt0rWsPckMNjKitP13nwC [0:3]; wire [16:0] Geu8JB9GQPz2V3cm3LHyYE [0:3]; wire Kkuw0xaU1gxu6c3MMwwn1E; wire signed [15:0] q1QqHpJturuPqVu8I4MkMSH; wire signed [15:0] q1WKxJkpU1brIIPGyF8fIVE; wire signed [15:0] iv8gJY2B57qsdytxw9VxiG; wire signed [15:0] lEFqYoOkSWU4q10gSVmI4E; wire signed [15:0] vMu9skGPdYyiM3oFdue24F; wire signed [15:0] xwezR2RIHC4PeBNYfGGfkC; wire signed [15:0] ULrCkIyU4pJmNi7CrWtDeF; wire signed [15:0] U4UeUPQOYvb97BDAB1FwND; wire signed [15:0] vVb1Nr8Z9IbM7qE1hxGtz [0:3]; wire signed [15:0] YFtm2iylQsm653bK0Hk0jH [0:3]; wire signed [15:0] Tr7iLo0EAESL4xlkesaUAF [0:3]; wire signed [15:0] p0O7euHBdo0osOt01nZPwG [0:3]; wire signed [15:0] JfSYs6vgqp2A4gS4D1psE; wire signed [15:0] iTlAzbO5ZYBZpOm5zhY7QG; wire signed [15:0] K5SwykB0asun0pcOcUmmXH; wire signed [15:0] IaiPYP7955Df4uWpAdYAzB; wire signed [15:0] b5TESZ6GeKtar9Blb1lj3OC; wire signed [15:0] v4tJvHK46bS3jIEwGDLaqnB; wire signed [15:0] eXq5fUFTZbAxieLoC9CpF; wire signed [15:0] d2SSAVXKXXa1w1k75YqDUH; wire signed [15:0] Sg3GG7AJ6DTTRqbnMxAozB [0:3]; wire signed [15:0] yUtorokxTduMdJFfTXXhnE [0:3]; wire k5IFxM0f5IPLItpTOfGOMG; wire signed [15:0] EIYK1nT0oJLxbcxjmodwrC; wire signed [15:0] l45qCeMpWMHOXjwYLaHORRE; wire signed [15:0] j8SzfGJHmeoXnV9bhAUk40F; wire signed [15:0] dMKGmQc7XAB1i3kk2Yk0hH; wire signed [15:0] ydI2XfENb2Kl0A3qJMSMBB; wire signed [15:0] nXMdpgmOgBwUAR30aQsd0B; wire signed [15:0] kenMGol9N3qu644VwSIQzD; wire signed [15:0] ovgS7leqdS5z2NH8xqTyeH; wire IwgDKbj92A15RKEkOdpXgE; reg [0:17] Fk3evzNcklSugbL51Yj8N; wire [0:17] k25NwHb1uJjT7flGGxsxBC; wire a2BLSsheDEDArqcNugKUoB; wire signed [15:0] ds3UaO1QhyfiWT7RZKX23G [0:3]; wire signed [15:0] tCCvu1nsVn6k0oKnEbNi9E [0:3]; wire [15:0] Vc8f45Qo75ucTzy0jKolzE; wire [15:0] ZNDiypKqoG4e82nJIljMu; wire [15:0] EW7O02E0JPjfI2XYnqHBZB; wire [15:0] b5ag7OG9oPVwNLOghEh9at; wire [15:0] rQqvnPiwzKpGmREAhe0vF [0:3]; wire cuj63SB5UdTmsBtbC9kwQH; wtU1sSRiRHqGwLWK3NzQmD mkKISPEnzvNlbXRBTQ83YC (.v04pHKxyc2sPW047bbyUgE(mclk), .JAMOfrNHxGSYDF0urqkLN(rstb), .r3faKvvHpwNbS8m4h6rXSUB(qdin_0), .cmM018LKGhcOIt4F15GJS(qdin_1), .J5kDQbkAAS4E39jPz9JzwD(qdin_2), .PVNB5uj77jMa2DXz4vJtIH(qdin_3), .xj2txhdk3kH1ioK0rKOVrG(f1en), .R6zf5iqRNVEGVBO8egq8kF(srst), .mdal5obekPJm0ao7ZiZ4cF(RDoofzNe0oXjNKPxTYnsJG), .q4mhS1P9mOTwehAXXNmhxF(l96ToZvA3JxZRoamoFQ1UB), .vyWRmDyKy2RVVIdRBtzV5F(vuBZeR1bCIQ7eYub4Nym0B), .SRoFC9yIIwEIUwYpoyy0QF(kYezVXe7e7E7TbchXde4QG), .wpHiLzmis5ns3l38MddOzE(BdTGl8ppsd8fNRyihNQvWD), .j963sPBld8mpm71sqcvb8WF(j5vaJTpXoIQ2WMB1cDQvqC), .Ic4vfYy6jnxaw8uXI98INH(fijzTATvD4NCVDjSoyqDXC), .x2KkW4HKTQgVBmVskDu4RD(uH5IsuPlvOkkvGQhI40ZZF), .g1D8wSsV4Ksuy5G0qxKYMs(TciTCDpCygk823aRzOkhCE) ); always @(posedge mclk or negedge rstb) begin : MJlo6U2223vRHOqbaXT3SB if (rstb == 1'b0) begin lYL40DZJNrZGA50HVltAXD <= 22'b0000000000000000000000; end else begin if (TciTCDpCygk823aRzOkhCE == 1'b1) begin if (lYL40DZJNrZGA50HVltAXD >= 22'b0001000000000000000000) begin lYL40DZJNrZGA50HVltAXD <= 22'b0000000000000000000000; end else begin lYL40DZJNrZGA50HVltAXD <= lYL40DZJNrZGA50HVltAXD + 22'b0000000000000000000001; end end end end assign d5CXluM5YmRNluM6LdzEuRD = {1'b0, {lYL40DZJNrZGA50HVltAXD, 21'b000000000000000000000}}; assign jAqDYspp5RSupfEc9vWoJH = d5CXluM5YmRNluM6LdzEuRD[36:19]; assign HHiAQq0eXS4V724AeWtEMD = jAqDYspp5RSupfEc9vWoJH >= 18'b100000000000000000; assign PFHmZS0ipZLKqJ39A27L8F = jAqDYspp5RSupfEc9vWoJH[16:0]; assign HtkwvAWd5V10OAKRmUTiLD = {15'b0, PFHmZS0ipZLKqJ39A27L8F}; assign IMy6yN0h9YqHeUl7378ZhB = HtkwvAWd5V10OAKRmUTiLD + 32'b00000000000000000000000000000011; assign FBdqgz94a8SGX1FULhpnhF = {1'b0, {IMy6yN0h9YqHeUl7378ZhB, 31'b0000000000000000000000000000000}}; assign eq6ExCvRAypD8ZXX1hJg2G = FBdqgz94a8SGX1FULhpnhF[50:41]; assign M6DCmjjEAXTHH63S0PcE0E = {22'b0, eq6ExCvRAypD8ZXX1hJg2G}; k67zvJy02k7XHYhPp3qIYH lH0t48igjoCV3d4v6rXTpC (.yQNwAzareGOhTeFAcGgFWE(M6DCmjjEAXTHH63S0PcE0E), .jqBlsvEQIekR8Gt2pzz5n(ImRl6qg5Qleo28k6kzf5ID) ); assign xWllAgKkXsJdEckAS1JkRE = {1'b0, {ImRl6qg5Qleo28k6kzf5ID, 15'b000000000000000}}; assign txIZVPOqyNjR0XJaNnEWgC = {6'b0, xWllAgKkXsJdEckAS1JkRE[31:21]}; assign o8JfccMcxN3IkRA878Wl6qB[0] = 17'b00000000000000011; assign o8JfccMcxN3IkRA878Wl6qB[1] = 17'b00000000000000010; assign o8JfccMcxN3IkRA878Wl6qB[2] = 17'b00000000000000001; assign o8JfccMcxN3IkRA878Wl6qB[3] = 17'b00000000000000000; assign iVUCRzTzoib1t9JQL19F1B[0] = txIZVPOqyNjR0XJaNnEWgC + o8JfccMcxN3IkRA878Wl6qB[0]; assign iVUCRzTzoib1t9JQL19F1B[1] = txIZVPOqyNjR0XJaNnEWgC + o8JfccMcxN3IkRA878Wl6qB[1]; assign iVUCRzTzoib1t9JQL19F1B[2] = txIZVPOqyNjR0XJaNnEWgC + o8JfccMcxN3IkRA878Wl6qB[2]; assign iVUCRzTzoib1t9JQL19F1B[3] = txIZVPOqyNjR0XJaNnEWgC + o8JfccMcxN3IkRA878Wl6qB[3]; assign q8UubaExFIU37MrHaKCYjEH[0] = iVUCRzTzoib1t9JQL19F1B[0][1:0]; assign q8UubaExFIU37MrHaKCYjEH[1] = iVUCRzTzoib1t9JQL19F1B[1][1:0]; assign q8UubaExFIU37MrHaKCYjEH[2] = iVUCRzTzoib1t9JQL19F1B[2][1:0]; assign q8UubaExFIU37MrHaKCYjEH[3] = iVUCRzTzoib1t9JQL19F1B[3][1:0]; assign i3T8rgFVbtYhLp11xyNVaG = {31'b0, q8UubaExFIU37MrHaKCYjEH[0]}; assign kmQDARJ5RSC33fkFkFEZvB[0] = 33'sh000000003 - i3T8rgFVbtYhLp11xyNVaG; assign xb5OWtSspXT5QIrsjYRNyC = {31'b0, q8UubaExFIU37MrHaKCYjEH[1]}; assign kmQDARJ5RSC33fkFkFEZvB[1] = 33'sh000000003 - xb5OWtSspXT5QIrsjYRNyC; assign zkeZd8GIm1z3m743ZzXwoF = {31'b0, q8UubaExFIU37MrHaKCYjEH[2]}; assign kmQDARJ5RSC33fkFkFEZvB[2] = 33'sh000000003 - zkeZd8GIm1z3m743ZzXwoF; assign d3io0lXPWPHhxjlWak3S1G = {31'b0, q8UubaExFIU37MrHaKCYjEH[3]}; assign kmQDARJ5RSC33fkFkFEZvB[3] = 33'sh000000003 - d3io0lXPWPHhxjlWak3S1G; assign h6X6Ift6lj74yXs2DyR91PG = {1'b0, {IMy6yN0h9YqHeUl7378ZhB, 31'b0000000000000000000000000000000}}; assign v0ZPFDd9cyRidUk0uUpeZF = {6'b0, h6X6Ift6lj74yXs2DyR91PG[63:38]}; e8HeF7GSPxfrhisMVdBBvN zqR2DjED1zsOu7YhFxEFnE (.yQNwAzareGOhTeFAcGgFWE(v0ZPFDd9cyRidUk0uUpeZF), .jqBlsvEQIekR8Gt2pzz5n(UGX8fdfHPAfRuWbIXSAJkC) ); assign iUgDeFg7wK7VmcsUejECJE = {1'b0, {UGX8fdfHPAfRuWbIXSAJkC, 15'b000000000000000}}; assign kXQPeGN2PPqOhoBeXJau8E = {3'b0, iUgDeFg7wK7VmcsUejECJE[31:18]}; assign RgAX8O9DbR6HNMiXsFyzb[0] = 17'b00000000000000000; assign RgAX8O9DbR6HNMiXsFyzb[1] = 17'b00000000000000001; assign RgAX8O9DbR6HNMiXsFyzb[2] = 17'b00000000000000010; assign RgAX8O9DbR6HNMiXsFyzb[3] = 17'b00000000000000011; assign Hm89BMHiz5dcKMTSyT6ZgE[0] = kXQPeGN2PPqOhoBeXJau8E + RgAX8O9DbR6HNMiXsFyzb[0]; assign Hm89BMHiz5dcKMTSyT6ZgE[1] = kXQPeGN2PPqOhoBeXJau8E + RgAX8O9DbR6HNMiXsFyzb[1]; assign Hm89BMHiz5dcKMTSyT6ZgE[2] = kXQPeGN2PPqOhoBeXJau8E + RgAX8O9DbR6HNMiXsFyzb[2]; assign Hm89BMHiz5dcKMTSyT6ZgE[3] = kXQPeGN2PPqOhoBeXJau8E + RgAX8O9DbR6HNMiXsFyzb[3]; assign TqEdytxeoETbv4LqQENvdE[0] = Hm89BMHiz5dcKMTSyT6ZgE[0][1:0]; assign TqEdytxeoETbv4LqQENvdE[1] = Hm89BMHiz5dcKMTSyT6ZgE[1][1:0]; assign TqEdytxeoETbv4LqQENvdE[2] = Hm89BMHiz5dcKMTSyT6ZgE[2][1:0]; assign TqEdytxeoETbv4LqQENvdE[3] = Hm89BMHiz5dcKMTSyT6ZgE[3][1:0]; assign HWvpOqHBtG8nHbtWWOs5ME[0] = {31'b0, TqEdytxeoETbv4LqQENvdE[0]}; assign HWvpOqHBtG8nHbtWWOs5ME[1] = {31'b0, TqEdytxeoETbv4LqQENvdE[1]}; assign HWvpOqHBtG8nHbtWWOs5ME[2] = {31'b0, TqEdytxeoETbv4LqQENvdE[2]}; assign HWvpOqHBtG8nHbtWWOs5ME[3] = {31'b0, TqEdytxeoETbv4LqQENvdE[3]}; assign XFDR6Vjpsj8y8if8sCJpyC[0] = (HHiAQq0eXS4V724AeWtEMD == 1'b0 ? kmQDARJ5RSC33fkFkFEZvB[0] : HWvpOqHBtG8nHbtWWOs5ME[0]); assign XFDR6Vjpsj8y8if8sCJpyC[1] = (HHiAQq0eXS4V724AeWtEMD == 1'b0 ? kmQDARJ5RSC33fkFkFEZvB[1] : HWvpOqHBtG8nHbtWWOs5ME[1]); assign XFDR6Vjpsj8y8if8sCJpyC[2] = (HHiAQq0eXS4V724AeWtEMD == 1'b0 ? kmQDARJ5RSC33fkFkFEZvB[2] : HWvpOqHBtG8nHbtWWOs5ME[2]); assign XFDR6Vjpsj8y8if8sCJpyC[3] = (HHiAQq0eXS4V724AeWtEMD == 1'b0 ? kmQDARJ5RSC33fkFkFEZvB[3] : HWvpOqHBtG8nHbtWWOs5ME[3]); always @(posedge mclk or negedge rstb) begin : b4269YDGE0N1rr5kDbvv4MG if (rstb == 1'b0) begin ZIXwDtDHOFCY284ItMUkPE[0] <= 33'sh000000000; ZIXwDtDHOFCY284ItMUkPE[1] <= 33'sh000000000; ZIXwDtDHOFCY284ItMUkPE[2] <= 33'sh000000000; ZIXwDtDHOFCY284ItMUkPE[3] <= 33'sh000000000; end else begin ZIXwDtDHOFCY284ItMUkPE[0] <= XFDR6Vjpsj8y8if8sCJpyC[0]; ZIXwDtDHOFCY284ItMUkPE[1] <= XFDR6Vjpsj8y8if8sCJpyC[1]; ZIXwDtDHOFCY284ItMUkPE[2] <= XFDR6Vjpsj8y8if8sCJpyC[2]; ZIXwDtDHOFCY284ItMUkPE[3] <= XFDR6Vjpsj8y8if8sCJpyC[3]; end end always @(posedge mclk or negedge rstb) begin : BI74HgUgswjF55jlBypAZE if (rstb == 1'b0) begin wmHZAgpaaD0AnBPdMzFAWB <= 1'b0; end else begin wmHZAgpaaD0AnBPdMzFAWB <= HHiAQq0eXS4V724AeWtEMD; end end assign JM1PWrdw4CsiaxhIFEj0FG[0] = PFHmZS0ipZLKqJ39A27L8F; assign JM1PWrdw4CsiaxhIFEj0FG[1] = PFHmZS0ipZLKqJ39A27L8F; assign JM1PWrdw4CsiaxhIFEj0FG[2] = PFHmZS0ipZLKqJ39A27L8F; assign JM1PWrdw4CsiaxhIFEj0FG[3] = PFHmZS0ipZLKqJ39A27L8F; assign NtsaMyVZXVYmztcjOvOk8 = {1'b0, {JM1PWrdw4CsiaxhIFEj0FG[0], 16'b0000000000000000}}; assign Bx5GbZBMMZWJmhJNe1plNE[0] = {1'b0, NtsaMyVZXVYmztcjOvOk8[33:18]}; assign Ow2gCZKYLWzsXB6jHnoqfG = {1'b0, {JM1PWrdw4CsiaxhIFEj0FG[1], 16'b0000000000000000}}; assign Bx5GbZBMMZWJmhJNe1plNE[1] = {1'b0, Ow2gCZKYLWzsXB6jHnoqfG[33:18]}; assign otv4IxbTPpKKTvscHxftHG = {1'b0, {JM1PWrdw4CsiaxhIFEj0FG[2], 16'b0000000000000000}}; assign Bx5GbZBMMZWJmhJNe1plNE[2] = {1'b0, otv4IxbTPpKKTvscHxftHG[33:18]}; assign l0guWc0JIHa1f8SBb77OlIC = {1'b0, {JM1PWrdw4CsiaxhIFEj0FG[3], 16'b0000000000000000}}; assign Bx5GbZBMMZWJmhJNe1plNE[3] = {1'b0, l0guWc0JIHa1f8SBb77OlIC[33:18]}; assign vDf5jyCbwqHvGEEIH52rqG[0] = {1'b0, Bx5GbZBMMZWJmhJNe1plNE[0]}; assign vDf5jyCbwqHvGEEIH52rqG[1] = {1'b0, Bx5GbZBMMZWJmhJNe1plNE[1]}; assign vDf5jyCbwqHvGEEIH52rqG[2] = {1'b0, Bx5GbZBMMZWJmhJNe1plNE[2]}; assign vDf5jyCbwqHvGEEIH52rqG[3] = {1'b0, Bx5GbZBMMZWJmhJNe1plNE[3]}; assign KyXrE6JYq7NUB9MlwmKcGH = HtkwvAWd5V10OAKRmUTiLD; assign THQEaifSmIkcouXcNP6X2G = HtkwvAWd5V10OAKRmUTiLD + 32'b00000000000000000000000000000001; assign Xp7jYGB4wGPVX0g6nIaYOD = HtkwvAWd5V10OAKRmUTiLD + 32'b00000000000000000000000000000010; xbcMJDB8htpX3R9YnKkaXC u3lZIgQMvq8uWQ6X01pbQ (.QQYO9noW2AzWAhLJIl3WIE(KyXrE6JYq7NUB9MlwmKcGH), .LIf9KkhuVKSu7vlUpWufBG(THQEaifSmIkcouXcNP6X2G), .c9WUZlfywHR3RaGJnbumYHB(Xp7jYGB4wGPVX0g6nIaYOD), .iU3uCiDXuU6z4nkTQ5PufE(IMy6yN0h9YqHeUl7378ZhB), .z8dRITT2PceChhB9z9EWBC(x2T5MHXEjHB4mbeunlQ5xlC), .N7ZKCQ4vfkUB2KkHwgE4GC(m3srRE1KQDnmVOjclDlFnB), .PfPBxRXyGunZRp8BSw7dcF(cZMBbP0tbfriJB96bWdXBG), .o5kjnQ9W5HT05kz0swOA6QH(OlmksAU0OqEmB1eHPlD4LF) ); assign wZQ5Nh8v8jyFGZaqm7MPFF[0] = x2T5MHXEjHB4mbeunlQ5xlC; assign wZQ5Nh8v8jyFGZaqm7MPFF[1] = m3srRE1KQDnmVOjclDlFnB; assign wZQ5Nh8v8jyFGZaqm7MPFF[2] = cZMBbP0tbfriJB96bWdXBG; assign wZQ5Nh8v8jyFGZaqm7MPFF[3] = OlmksAU0OqEmB1eHPlD4LF; assign K2KmCTF5G7ost89y9oqLiD = {1'b0, {wZQ5Nh8v8jyFGZaqm7MPFF[0], 15'b000000000000000}}; assign n7lC0EX54a5Db2Ey78BZWH[0] = {3'b0, K2KmCTF5G7ost89y9oqLiD[31:18]}; assign AIcGcubjt3yRVo2TP54CyG = {1'b0, {wZQ5Nh8v8jyFGZaqm7MPFF[1], 15'b000000000000000}}; assign n7lC0EX54a5Db2Ey78BZWH[1] = {3'b0, AIcGcubjt3yRVo2TP54CyG[31:18]}; assign DPfpo6Ze4IPKLEjjyJWtJD = {1'b0, {wZQ5Nh8v8jyFGZaqm7MPFF[2], 15'b000000000000000}}; assign n7lC0EX54a5Db2Ey78BZWH[2] = {3'b0, DPfpo6Ze4IPKLEjjyJWtJD[31:18]}; assign DKFv0pTB8YURDrEOItHrZH = {1'b0, {wZQ5Nh8v8jyFGZaqm7MPFF[3], 15'b000000000000000}}; assign n7lC0EX54a5Db2Ey78BZWH[3] = {3'b0, DKFv0pTB8YURDrEOItHrZH[31:18]}; assign gjjq7XRjRpkPoRKYu5l6n = {1'b0, {n7lC0EX54a5Db2Ey78BZWH[0], 16'b0000000000000000}}; assign mhinOy8fRr1hyDeV9qCPFB[0] = gjjq7XRjRpkPoRKYu5l6n[27:11]; assign hvpZkEPsH8kWqLanUTpxMB = {1'b0, {n7lC0EX54a5Db2Ey78BZWH[1], 16'b0000000000000000}}; assign mhinOy8fRr1hyDeV9qCPFB[1] = hvpZkEPsH8kWqLanUTpxMB[27:11]; assign zmbkHL82PolXRAHTmnIS9D = {1'b0, {n7lC0EX54a5Db2Ey78BZWH[2], 16'b0000000000000000}}; assign mhinOy8fRr1hyDeV9qCPFB[2] = zmbkHL82PolXRAHTmnIS9D[27:11]; assign g9yIixLFTxnivPa0KqVeY1D = {1'b0, {n7lC0EX54a5Db2Ey78BZWH[3], 16'b0000000000000000}}; assign mhinOy8fRr1hyDeV9qCPFB[3] = g9yIixLFTxnivPa0KqVeY1D[27:11]; assign ATVtgjciSvCRUI7H3Y9tuD = {1'b0, {txIZVPOqyNjR0XJaNnEWgC, 16'b0000000000000000}}; assign toucxMaGXtuei4mJhB7SvH = ATVtgjciSvCRUI7H3Y9tuD[27:18]; assign t1mfqjXjUa0cnuylRz3bBNF = {8'b0, toucxMaGXtuei4mJhB7SvH}; assign BQWUnHpxPEGrMvfoEg50BE[0] = ({1'b0, mhinOy8fRr1hyDeV9qCPFB[0]}) + t1mfqjXjUa0cnuylRz3bBNF; assign BQWUnHpxPEGrMvfoEg50BE[1] = ({1'b0, mhinOy8fRr1hyDeV9qCPFB[1]}) + t1mfqjXjUa0cnuylRz3bBNF; assign BQWUnHpxPEGrMvfoEg50BE[2] = ({1'b0, mhinOy8fRr1hyDeV9qCPFB[2]}) + t1mfqjXjUa0cnuylRz3bBNF; assign BQWUnHpxPEGrMvfoEg50BE[3] = ({1'b0, mhinOy8fRr1hyDeV9qCPFB[3]}) + t1mfqjXjUa0cnuylRz3bBNF; UoUhxjuVDf73mwAaAcjVRH JYlyLmYe4aXPfUjLR66lvF (.tu9ohhJdK00us7wfvWNQYC(XFDR6Vjpsj8y8if8sCJpyC[0]), .utKZyKAnyhCUOZ6LUagX4D(XFDR6Vjpsj8y8if8sCJpyC[1]), .gA7z08sAKJH0Dq3fae8ZeF(XFDR6Vjpsj8y8if8sCJpyC[2]), .vrNoBb2ZnRj9xKaojUq7EG(XFDR6Vjpsj8y8if8sCJpyC[3]), .b0y2UtjO5W56S6DbL4mEOC(BQWUnHpxPEGrMvfoEg50BE[0]), .Htw4jhVkz8IRnd9IbKpIUC(BQWUnHpxPEGrMvfoEg50BE[1]), .y4o9opauBD4PXZzgZLUETHF(BQWUnHpxPEGrMvfoEg50BE[2]), .yPz5e3igECVkjPPXSkoiHG(BQWUnHpxPEGrMvfoEg50BE[3]), .z8dRITT2PceChhB9z9EWBC(UIikZeafI7JRbAIwWZXxZG), .N7ZKCQ4vfkUB2KkHwgE4GC(YHsZm9RxIvVHFFCFqjHJbB), .PfPBxRXyGunZRp8BSw7dcF(Ro8Qq6Y03XDjqsnyirVcTD), .o5kjnQ9W5HT05kz0swOA6QH(XW2XizJGnQkUYhMVZ7vzD) ); assign KRGfxNqFr6P3qLzrH4DIYD[0] = UIikZeafI7JRbAIwWZXxZG; assign KRGfxNqFr6P3qLzrH4DIYD[1] = YHsZm9RxIvVHFFCFqjHJbB; assign KRGfxNqFr6P3qLzrH4DIYD[2] = Ro8Qq6Y03XDjqsnyirVcTD; assign KRGfxNqFr6P3qLzrH4DIYD[3] = XW2XizJGnQkUYhMVZ7vzD; assign YkB06NLyXnKPFxzf13DnpH[0] = (HHiAQq0eXS4V724AeWtEMD == 1'b0 ? vDf5jyCbwqHvGEEIH52rqG[0] : KRGfxNqFr6P3qLzrH4DIYD[0]); assign YkB06NLyXnKPFxzf13DnpH[1] = (HHiAQq0eXS4V724AeWtEMD == 1'b0 ? vDf5jyCbwqHvGEEIH52rqG[1] : KRGfxNqFr6P3qLzrH4DIYD[1]); assign YkB06NLyXnKPFxzf13DnpH[2] = (HHiAQq0eXS4V724AeWtEMD == 1'b0 ? vDf5jyCbwqHvGEEIH52rqG[2] : KRGfxNqFr6P3qLzrH4DIYD[2]); assign YkB06NLyXnKPFxzf13DnpH[3] = (HHiAQq0eXS4V724AeWtEMD == 1'b0 ? vDf5jyCbwqHvGEEIH52rqG[3] : KRGfxNqFr6P3qLzrH4DIYD[3]); assign gAw9zJNNZqPQfnlAoc3jXH[0] = YkB06NLyXnKPFxzf13DnpH[0][16:0]; assign gAw9zJNNZqPQfnlAoc3jXH[1] = YkB06NLyXnKPFxzf13DnpH[1][16:0]; assign gAw9zJNNZqPQfnlAoc3jXH[2] = YkB06NLyXnKPFxzf13DnpH[2][16:0]; assign gAw9zJNNZqPQfnlAoc3jXH[3] = YkB06NLyXnKPFxzf13DnpH[3][16:0]; assign CqX3zbRXkD0JZjUDCE4uyC[0] = RDoofzNe0oXjNKPxTYnsJG; assign CqX3zbRXkD0JZjUDCE4uyC[1] = l96ToZvA3JxZRoamoFQ1UB; assign CqX3zbRXkD0JZjUDCE4uyC[2] = vuBZeR1bCIQ7eYub4Nym0B; assign CqX3zbRXkD0JZjUDCE4uyC[3] = kYezVXe7e7E7TbchXde4QG; assign Y2qRC0lD6WkLUd7tO2DL8D[0] = BdTGl8ppsd8fNRyihNQvWD; assign Y2qRC0lD6WkLUd7tO2DL8D[1] = j5vaJTpXoIQ2WMB1cDQvqC; assign Y2qRC0lD6WkLUd7tO2DL8D[2] = fijzTATvD4NCVDjSoyqDXC; assign Y2qRC0lD6WkLUd7tO2DL8D[3] = uH5IsuPlvOkkvGQhI40ZZF; n0XvT1ntWfPOHFF4mUMwzZ pxchbFl1AiSqRZyg96cup (.tu9ohhJdK00us7wfvWNQYC(XFDR6Vjpsj8y8if8sCJpyC[0]), .utKZyKAnyhCUOZ6LUagX4D(XFDR6Vjpsj8y8if8sCJpyC[1]), .gA7z08sAKJH0Dq3fae8ZeF(XFDR6Vjpsj8y8if8sCJpyC[2]), .vrNoBb2ZnRj9xKaojUq7EG(XFDR6Vjpsj8y8if8sCJpyC[3]), .IS0z2hJ2LtWljhJ4YYLYaE(CqX3zbRXkD0JZjUDCE4uyC[0]), .TkIATgh1a29iglca8RarC(CqX3zbRXkD0JZjUDCE4uyC[1]), .b4TwkCZxxInAgelXDhMy8E(CqX3zbRXkD0JZjUDCE4uyC[2]), .f9IpN1esn9PJkU40eAffHB(CqX3zbRXkD0JZjUDCE4uyC[3]), .ySOrNaQmYucOX4cyOT5LnG(Y2qRC0lD6WkLUd7tO2DL8D[0]), .gmoWrkWFJMiyePfRw5V1lD(Y2qRC0lD6WkLUd7tO2DL8D[1]), .nzbLrBOekdX928cLtCU5jD(Y2qRC0lD6WkLUd7tO2DL8D[2]), .a9DSedGWFdieeZlu7mhtF7D(Y2qRC0lD6WkLUd7tO2DL8D[3]), .zzBKVZ6VX4ht5u9x9EjCiD(w27urwsxsx3vX1J4eEaqy0D), .j83GXtGY1eMU252JJ6B9mC(onEIj0VH5ehJOImYn9CHFC), .r7Q5mFJeRMLiOPMHQDcQQB(GyXnWgCHVjevCAC5dsEk8G), .wtshVXYU5akP8bsJW8meZH(dCpVrDZOfokUK9iu0jbwzC), .w2g8aZ7DNLiB7xd9ema9tID(h8Njhoqboql6ktvl74YNlD), .EpypH5ZIz8rvw2qkajrEUD(g0CmNQp5HtaKwsfnggkLOD), .k5yT5mPpUVKMKN3fkRm1LR(r7YnXgwRbNGWdEl2TZcAw0C), .hfxEgMPHtdNs5za4aJfZR(u1xFlD3D83sqzZNknRicP6B) ); kkELk45BoVareqHanLSiwD NFIAvWAmRi26bAmV4HqixB (.rstb(rstb), .v04pHKxyc2sPW047bbyUgE(mclk), .vLtlRIKgN8j1pwmLLNsPG(gAw9zJNNZqPQfnlAoc3jXH[0]), .JzMAX1dysSuDOcRjDKM6jE(gAw9zJNNZqPQfnlAoc3jXH[1]), .mFPagULjpfgerkfoXcLj6E(gAw9zJNNZqPQfnlAoc3jXH[2]), .ZxXeSJVdqJaLdxkVQHDcKE(gAw9zJNNZqPQfnlAoc3jXH[3]), .m5wgqFuUcW1FOMsh4Ru6H(w27urwsxsx3vX1J4eEaqy0D), .KMtac8skVU06MkqFCILXMF(onEIj0VH5ehJOImYn9CHFC), .n3sKmw6MRNFgYu3FVurx4gF(GyXnWgCHVjevCAC5dsEk8G), .ruH3uKgP1LYhGZv6tkbvYB(dCpVrDZOfokUK9iu0jbwzC), .h5UJTRfxlrAz6m3sECIknXE(h8Njhoqboql6ktvl74YNlD), .Fr5Lz9pdsoRhxTCNFip6AE(g0CmNQp5HtaKwsfnggkLOD), .uG1VLsSqDTRiixegby6clE(r7YnXgwRbNGWdEl2TZcAw0C), .qqi4ViVQH4ZOVdWVypt4yB(u1xFlD3D83sqzZNknRicP6B), .UKo8akspo4h0jsZ6g712NB(HHiAQq0eXS4V724AeWtEMD), .zzBKVZ6VX4ht5u9x9EjCiD(M5pFttxc4QndsuSd89rKrD), .j83GXtGY1eMU252JJ6B9mC(FVvSvaFiVsOXZzGo86bsoC), .r7Q5mFJeRMLiOPMHQDcQQB(dte5acyHW51RNSwjPM8XJD), .wtshVXYU5akP8bsJW8meZH(wLogEYXttTcYn1hYyKkIwE), .w2g8aZ7DNLiB7xd9ema9tID(Z1XJpcLo4zUnViPcNLmlmC), .EpypH5ZIz8rvw2qkajrEUD(yfb14sul5mbLBMqiwceCCC), .k5yT5mPpUVKMKN3fkRm1LR(nz8qYIrRTZKfZJZAE7BZrF), .hfxEgMPHtdNs5za4aJfZR(iZEHwpNoTE4xYjGNgFVDSH) ); assign AvHKfOLcDBK6tGfufEsPhF[0] = M5pFttxc4QndsuSd89rKrD; assign AvHKfOLcDBK6tGfufEsPhF[1] = FVvSvaFiVsOXZzGo86bsoC; assign AvHKfOLcDBK6tGfufEsPhF[2] = dte5acyHW51RNSwjPM8XJD; assign AvHKfOLcDBK6tGfufEsPhF[3] = wLogEYXttTcYn1hYyKkIwE; assign AUkBI5w4Pfinl5l6Ts0oXB[0] = Z1XJpcLo4zUnViPcNLmlmC; assign AUkBI5w4Pfinl5l6Ts0oXB[1] = yfb14sul5mbLBMqiwceCCC; assign AUkBI5w4Pfinl5l6Ts0oXB[2] = nz8qYIrRTZKfZJZAE7BZrF; assign AUkBI5w4Pfinl5l6Ts0oXB[3] = iZEHwpNoTE4xYjGNgFVDSH; assign perQtgyUzTQmgJPDhQgq5D[0] = {1'b0, Bx5GbZBMMZWJmhJNe1plNE[0]}; assign perQtgyUzTQmgJPDhQgq5D[1] = {1'b0, Bx5GbZBMMZWJmhJNe1plNE[1]}; assign perQtgyUzTQmgJPDhQgq5D[2] = {1'b0, Bx5GbZBMMZWJmhJNe1plNE[2]}; assign perQtgyUzTQmgJPDhQgq5D[3] = {1'b0, Bx5GbZBMMZWJmhJNe1plNE[3]}; assign wnt0rWsPckMNjKitP13nwC[0] = (HHiAQq0eXS4V724AeWtEMD == 1'b0 ? KRGfxNqFr6P3qLzrH4DIYD[0] : perQtgyUzTQmgJPDhQgq5D[0]); assign wnt0rWsPckMNjKitP13nwC[1] = (HHiAQq0eXS4V724AeWtEMD == 1'b0 ? KRGfxNqFr6P3qLzrH4DIYD[1] : perQtgyUzTQmgJPDhQgq5D[1]); assign wnt0rWsPckMNjKitP13nwC[2] = (HHiAQq0eXS4V724AeWtEMD == 1'b0 ? KRGfxNqFr6P3qLzrH4DIYD[2] : perQtgyUzTQmgJPDhQgq5D[2]); assign wnt0rWsPckMNjKitP13nwC[3] = (HHiAQq0eXS4V724AeWtEMD == 1'b0 ? KRGfxNqFr6P3qLzrH4DIYD[3] : perQtgyUzTQmgJPDhQgq5D[3]); assign Geu8JB9GQPz2V3cm3LHyYE[0] = wnt0rWsPckMNjKitP13nwC[0][16:0]; assign Geu8JB9GQPz2V3cm3LHyYE[1] = wnt0rWsPckMNjKitP13nwC[1][16:0]; assign Geu8JB9GQPz2V3cm3LHyYE[2] = wnt0rWsPckMNjKitP13nwC[2][16:0]; assign Geu8JB9GQPz2V3cm3LHyYE[3] = wnt0rWsPckMNjKitP13nwC[3][16:0]; assign Kkuw0xaU1gxu6c3MMwwn1E = ~ HHiAQq0eXS4V724AeWtEMD; kkELk45BoVareqHanLSiwD Ymxl29V1ihNRAdK2DEWUhH (.rstb(rstb), .v04pHKxyc2sPW047bbyUgE(mclk), .vLtlRIKgN8j1pwmLLNsPG(Geu8JB9GQPz2V3cm3LHyYE[0]), .JzMAX1dysSuDOcRjDKM6jE(Geu8JB9GQPz2V3cm3LHyYE[1]), .mFPagULjpfgerkfoXcLj6E(Geu8JB9GQPz2V3cm3LHyYE[2]), .ZxXeSJVdqJaLdxkVQHDcKE(Geu8JB9GQPz2V3cm3LHyYE[3]), .m5wgqFuUcW1FOMsh4Ru6H(w27urwsxsx3vX1J4eEaqy0D), .KMtac8skVU06MkqFCILXMF(onEIj0VH5ehJOImYn9CHFC), .n3sKmw6MRNFgYu3FVurx4gF(GyXnWgCHVjevCAC5dsEk8G), .ruH3uKgP1LYhGZv6tkbvYB(dCpVrDZOfokUK9iu0jbwzC), .h5UJTRfxlrAz6m3sECIknXE(h8Njhoqboql6ktvl74YNlD), .Fr5Lz9pdsoRhxTCNFip6AE(g0CmNQp5HtaKwsfnggkLOD), .uG1VLsSqDTRiixegby6clE(r7YnXgwRbNGWdEl2TZcAw0C), .qqi4ViVQH4ZOVdWVypt4yB(u1xFlD3D83sqzZNknRicP6B), .UKo8akspo4h0jsZ6g712NB(Kkuw0xaU1gxu6c3MMwwn1E), .zzBKVZ6VX4ht5u9x9EjCiD(q1QqHpJturuPqVu8I4MkMSH), .j83GXtGY1eMU252JJ6B9mC(q1WKxJkpU1brIIPGyF8fIVE), .r7Q5mFJeRMLiOPMHQDcQQB(iv8gJY2B57qsdytxw9VxiG), .wtshVXYU5akP8bsJW8meZH(lEFqYoOkSWU4q10gSVmI4E), .w2g8aZ7DNLiB7xd9ema9tID(vMu9skGPdYyiM3oFdue24F), .EpypH5ZIz8rvw2qkajrEUD(xwezR2RIHC4PeBNYfGGfkC), .k5yT5mPpUVKMKN3fkRm1LR(ULrCkIyU4pJmNi7CrWtDeF), .hfxEgMPHtdNs5za4aJfZR(U4UeUPQOYvb97BDAB1FwND) ); assign vVb1Nr8Z9IbM7qE1hxGtz[0] = q1QqHpJturuPqVu8I4MkMSH; assign vVb1Nr8Z9IbM7qE1hxGtz[1] = q1WKxJkpU1brIIPGyF8fIVE; assign vVb1Nr8Z9IbM7qE1hxGtz[2] = iv8gJY2B57qsdytxw9VxiG; assign vVb1Nr8Z9IbM7qE1hxGtz[3] = lEFqYoOkSWU4q10gSVmI4E; assign YFtm2iylQsm653bK0Hk0jH[0] = vMu9skGPdYyiM3oFdue24F; assign YFtm2iylQsm653bK0Hk0jH[1] = xwezR2RIHC4PeBNYfGGfkC; assign YFtm2iylQsm653bK0Hk0jH[2] = ULrCkIyU4pJmNi7CrWtDeF; assign YFtm2iylQsm653bK0Hk0jH[3] = U4UeUPQOYvb97BDAB1FwND; assign Tr7iLo0EAESL4xlkesaUAF[0] = (wmHZAgpaaD0AnBPdMzFAWB == 1'b0 ? AvHKfOLcDBK6tGfufEsPhF[0] : vVb1Nr8Z9IbM7qE1hxGtz[0]); assign Tr7iLo0EAESL4xlkesaUAF[1] = (wmHZAgpaaD0AnBPdMzFAWB == 1'b0 ? AvHKfOLcDBK6tGfufEsPhF[1] : vVb1Nr8Z9IbM7qE1hxGtz[1]); assign Tr7iLo0EAESL4xlkesaUAF[2] = (wmHZAgpaaD0AnBPdMzFAWB == 1'b0 ? AvHKfOLcDBK6tGfufEsPhF[2] : vVb1Nr8Z9IbM7qE1hxGtz[2]); assign Tr7iLo0EAESL4xlkesaUAF[3] = (wmHZAgpaaD0AnBPdMzFAWB == 1'b0 ? AvHKfOLcDBK6tGfufEsPhF[3] : vVb1Nr8Z9IbM7qE1hxGtz[3]); assign p0O7euHBdo0osOt01nZPwG[0] = (wmHZAgpaaD0AnBPdMzFAWB == 1'b0 ? AUkBI5w4Pfinl5l6Ts0oXB[0] : YFtm2iylQsm653bK0Hk0jH[0]); assign p0O7euHBdo0osOt01nZPwG[1] = (wmHZAgpaaD0AnBPdMzFAWB == 1'b0 ? AUkBI5w4Pfinl5l6Ts0oXB[1] : YFtm2iylQsm653bK0Hk0jH[1]); assign p0O7euHBdo0osOt01nZPwG[2] = (wmHZAgpaaD0AnBPdMzFAWB == 1'b0 ? AUkBI5w4Pfinl5l6Ts0oXB[2] : YFtm2iylQsm653bK0Hk0jH[2]); assign p0O7euHBdo0osOt01nZPwG[3] = (wmHZAgpaaD0AnBPdMzFAWB == 1'b0 ? AUkBI5w4Pfinl5l6Ts0oXB[3] : YFtm2iylQsm653bK0Hk0jH[3]); QCP2KsVCXOv9pucMwLlsBG RW9qYuU77YZzJYTumStZh (.tu9ohhJdK00us7wfvWNQYC(ZIXwDtDHOFCY284ItMUkPE[0]), .utKZyKAnyhCUOZ6LUagX4D(ZIXwDtDHOFCY284ItMUkPE[1]), .gA7z08sAKJH0Dq3fae8ZeF(ZIXwDtDHOFCY284ItMUkPE[2]), .vrNoBb2ZnRj9xKaojUq7EG(ZIXwDtDHOFCY284ItMUkPE[3]), .IS0z2hJ2LtWljhJ4YYLYaE(Tr7iLo0EAESL4xlkesaUAF[0]), .TkIATgh1a29iglca8RarC(Tr7iLo0EAESL4xlkesaUAF[1]), .b4TwkCZxxInAgelXDhMy8E(Tr7iLo0EAESL4xlkesaUAF[2]), .f9IpN1esn9PJkU40eAffHB(Tr7iLo0EAESL4xlkesaUAF[3]), .ySOrNaQmYucOX4cyOT5LnG(p0O7euHBdo0osOt01nZPwG[0]), .gmoWrkWFJMiyePfRw5V1lD(p0O7euHBdo0osOt01nZPwG[1]), .nzbLrBOekdX928cLtCU5jD(p0O7euHBdo0osOt01nZPwG[2]), .a9DSedGWFdieeZlu7mhtF7D(p0O7euHBdo0osOt01nZPwG[3]), .zzBKVZ6VX4ht5u9x9EjCiD(JfSYs6vgqp2A4gS4D1psE), .j83GXtGY1eMU252JJ6B9mC(iTlAzbO5ZYBZpOm5zhY7QG), .r7Q5mFJeRMLiOPMHQDcQQB(K5SwykB0asun0pcOcUmmXH), .wtshVXYU5akP8bsJW8meZH(IaiPYP7955Df4uWpAdYAzB), .w2g8aZ7DNLiB7xd9ema9tID(b5TESZ6GeKtar9Blb1lj3OC), .EpypH5ZIz8rvw2qkajrEUD(v4tJvHK46bS3jIEwGDLaqnB), .k5yT5mPpUVKMKN3fkRm1LR(eXq5fUFTZbAxieLoC9CpF), .hfxEgMPHtdNs5za4aJfZR(d2SSAVXKXXa1w1k75YqDUH) ); assign Sg3GG7AJ6DTTRqbnMxAozB[0] = JfSYs6vgqp2A4gS4D1psE; assign Sg3GG7AJ6DTTRqbnMxAozB[1] = iTlAzbO5ZYBZpOm5zhY7QG; assign Sg3GG7AJ6DTTRqbnMxAozB[2] = K5SwykB0asun0pcOcUmmXH; assign Sg3GG7AJ6DTTRqbnMxAozB[3] = IaiPYP7955Df4uWpAdYAzB; assign yUtorokxTduMdJFfTXXhnE[0] = b5TESZ6GeKtar9Blb1lj3OC; assign yUtorokxTduMdJFfTXXhnE[1] = v4tJvHK46bS3jIEwGDLaqnB; assign yUtorokxTduMdJFfTXXhnE[2] = eXq5fUFTZbAxieLoC9CpF; assign yUtorokxTduMdJFfTXXhnE[3] = d2SSAVXKXXa1w1k75YqDUH; assign k5IFxM0f5IPLItpTOfGOMG = lYL40DZJNrZGA50HVltAXD >= 22'b0000001000000000000001; d4QD8esP7XdYbm4O3mpV7GH SeEGwQ0moTiTHYs4BaN8MC (.v04pHKxyc2sPW047bbyUgE(mclk), .JAMOfrNHxGSYDF0urqkLN(rstb), .w3gGIVls9UktX3B50XtCM9D(Sg3GG7AJ6DTTRqbnMxAozB[0]), .PkjFB7tzez7RAWc2cSLnBD(Sg3GG7AJ6DTTRqbnMxAozB[1]), .cuDt5zGIRdJYB1ZsmaWyNE(Sg3GG7AJ6DTTRqbnMxAozB[2]), .a1hhzPnRvmngQQ69MdICU7C(Sg3GG7AJ6DTTRqbnMxAozB[3]), .PF6wwTYP1q9nJ5YwMDlzXE(yUtorokxTduMdJFfTXXhnE[0]), .NunEp0PDJBOuCyVdY3ejIC(yUtorokxTduMdJFfTXXhnE[1]), .zTC5dHloAQWrunmpBf9AuG(yUtorokxTduMdJFfTXXhnE[2]), .d8pq1PMmLZANfmOanWWlBYF(yUtorokxTduMdJFfTXXhnE[3]), .xj2txhdk3kH1ioK0rKOVrG(k5IFxM0f5IPLItpTOfGOMG), .R6zf5iqRNVEGVBO8egq8kF(srst), .mdal5obekPJm0ao7ZiZ4cF(EIYK1nT0oJLxbcxjmodwrC), .q4mhS1P9mOTwehAXXNmhxF(l45qCeMpWMHOXjwYLaHORRE), .vyWRmDyKy2RVVIdRBtzV5F(j8SzfGJHmeoXnV9bhAUk40F), .SRoFC9yIIwEIUwYpoyy0QF(dMKGmQc7XAB1i3kk2Yk0hH), .wpHiLzmis5ns3l38MddOzE(ydI2XfENb2Kl0A3qJMSMBB), .j963sPBld8mpm71sqcvb8WF(nXMdpgmOgBwUAR30aQsd0B), .Ic4vfYy6jnxaw8uXI98INH(kenMGol9N3qu644VwSIQzD), .x2KkW4HKTQgVBmVskDu4RD(ovgS7leqdS5z2NH8xqTyeH), .g1D8wSsV4Ksuy5G0qxKYMs(IwgDKbj92A15RKEkOdpXgE) ); always @(posedge mclk or negedge rstb) begin : c4aO26E6Iq0zAPPqlEtwKoE if (rstb == 1'b0) begin Fk3evzNcklSugbL51Yj8N[0] <= 1'b0; Fk3evzNcklSugbL51Yj8N[1] <= 1'b0; Fk3evzNcklSugbL51Yj8N[2] <= 1'b0; Fk3evzNcklSugbL51Yj8N[3] <= 1'b0; Fk3evzNcklSugbL51Yj8N[4] <= 1'b0; Fk3evzNcklSugbL51Yj8N[5] <= 1'b0; Fk3evzNcklSugbL51Yj8N[6] <= 1'b0; Fk3evzNcklSugbL51Yj8N[7] <= 1'b0; Fk3evzNcklSugbL51Yj8N[8] <= 1'b0; Fk3evzNcklSugbL51Yj8N[9] <= 1'b0; Fk3evzNcklSugbL51Yj8N[10] <= 1'b0; Fk3evzNcklSugbL51Yj8N[11] <= 1'b0; Fk3evzNcklSugbL51Yj8N[12] <= 1'b0; Fk3evzNcklSugbL51Yj8N[13] <= 1'b0; Fk3evzNcklSugbL51Yj8N[14] <= 1'b0; Fk3evzNcklSugbL51Yj8N[15] <= 1'b0; Fk3evzNcklSugbL51Yj8N[16] <= 1'b0; Fk3evzNcklSugbL51Yj8N[17] <= 1'b0; end else begin Fk3evzNcklSugbL51Yj8N[0] <= k25NwHb1uJjT7flGGxsxBC[0]; Fk3evzNcklSugbL51Yj8N[1] <= k25NwHb1uJjT7flGGxsxBC[1]; Fk3evzNcklSugbL51Yj8N[2] <= k25NwHb1uJjT7flGGxsxBC[2]; Fk3evzNcklSugbL51Yj8N[3] <= k25NwHb1uJjT7flGGxsxBC[3]; Fk3evzNcklSugbL51Yj8N[4] <= k25NwHb1uJjT7flGGxsxBC[4]; Fk3evzNcklSugbL51Yj8N[5] <= k25NwHb1uJjT7flGGxsxBC[5]; Fk3evzNcklSugbL51Yj8N[6] <= k25NwHb1uJjT7flGGxsxBC[6]; Fk3evzNcklSugbL51Yj8N[7] <= k25NwHb1uJjT7flGGxsxBC[7]; Fk3evzNcklSugbL51Yj8N[8] <= k25NwHb1uJjT7flGGxsxBC[8]; Fk3evzNcklSugbL51Yj8N[9] <= k25NwHb1uJjT7flGGxsxBC[9]; Fk3evzNcklSugbL51Yj8N[10] <= k25NwHb1uJjT7flGGxsxBC[10]; Fk3evzNcklSugbL51Yj8N[11] <= k25NwHb1uJjT7flGGxsxBC[11]; Fk3evzNcklSugbL51Yj8N[12] <= k25NwHb1uJjT7flGGxsxBC[12]; Fk3evzNcklSugbL51Yj8N[13] <= k25NwHb1uJjT7flGGxsxBC[13]; Fk3evzNcklSugbL51Yj8N[14] <= k25NwHb1uJjT7flGGxsxBC[14]; Fk3evzNcklSugbL51Yj8N[15] <= k25NwHb1uJjT7flGGxsxBC[15]; Fk3evzNcklSugbL51Yj8N[16] <= k25NwHb1uJjT7flGGxsxBC[16]; Fk3evzNcklSugbL51Yj8N[17] <= k25NwHb1uJjT7flGGxsxBC[17]; end end assign a2BLSsheDEDArqcNugKUoB = Fk3evzNcklSugbL51Yj8N[17]; assign k25NwHb1uJjT7flGGxsxBC[0] = IwgDKbj92A15RKEkOdpXgE; assign k25NwHb1uJjT7flGGxsxBC[1] = Fk3evzNcklSugbL51Yj8N[0]; assign k25NwHb1uJjT7flGGxsxBC[2] = Fk3evzNcklSugbL51Yj8N[1]; assign k25NwHb1uJjT7flGGxsxBC[3] = Fk3evzNcklSugbL51Yj8N[2]; assign k25NwHb1uJjT7flGGxsxBC[4] = Fk3evzNcklSugbL51Yj8N[3]; assign k25NwHb1uJjT7flGGxsxBC[5] = Fk3evzNcklSugbL51Yj8N[4]; assign k25NwHb1uJjT7flGGxsxBC[6] = Fk3evzNcklSugbL51Yj8N[5]; assign k25NwHb1uJjT7flGGxsxBC[7] = Fk3evzNcklSugbL51Yj8N[6]; assign k25NwHb1uJjT7flGGxsxBC[8] = Fk3evzNcklSugbL51Yj8N[7]; assign k25NwHb1uJjT7flGGxsxBC[9] = Fk3evzNcklSugbL51Yj8N[8]; assign k25NwHb1uJjT7flGGxsxBC[10] = Fk3evzNcklSugbL51Yj8N[9]; assign k25NwHb1uJjT7flGGxsxBC[11] = Fk3evzNcklSugbL51Yj8N[10]; assign k25NwHb1uJjT7flGGxsxBC[12] = Fk3evzNcklSugbL51Yj8N[11]; assign k25NwHb1uJjT7flGGxsxBC[13] = Fk3evzNcklSugbL51Yj8N[12]; assign k25NwHb1uJjT7flGGxsxBC[14] = Fk3evzNcklSugbL51Yj8N[13]; assign k25NwHb1uJjT7flGGxsxBC[15] = Fk3evzNcklSugbL51Yj8N[14]; assign k25NwHb1uJjT7flGGxsxBC[16] = Fk3evzNcklSugbL51Yj8N[15]; assign k25NwHb1uJjT7flGGxsxBC[17] = Fk3evzNcklSugbL51Yj8N[16]; assign f2Vld = a2BLSsheDEDArqcNugKUoB; assign ds3UaO1QhyfiWT7RZKX23G[0] = EIYK1nT0oJLxbcxjmodwrC; assign ds3UaO1QhyfiWT7RZKX23G[1] = l45qCeMpWMHOXjwYLaHORRE; assign ds3UaO1QhyfiWT7RZKX23G[2] = j8SzfGJHmeoXnV9bhAUk40F; assign ds3UaO1QhyfiWT7RZKX23G[3] = dMKGmQc7XAB1i3kk2Yk0hH; assign tCCvu1nsVn6k0oKnEbNi9E[0] = ydI2XfENb2Kl0A3qJMSMBB; assign tCCvu1nsVn6k0oKnEbNi9E[1] = nXMdpgmOgBwUAR30aQsd0B; assign tCCvu1nsVn6k0oKnEbNi9E[2] = kenMGol9N3qu644VwSIQzD; assign tCCvu1nsVn6k0oKnEbNi9E[3] = ovgS7leqdS5z2NH8xqTyeH; yp36yVdBki2iBRVFYzbmt wctO69sGqqXIDGOi3l1nWB (.v04pHKxyc2sPW047bbyUgE(mclk), .JAMOfrNHxGSYDF0urqkLN(rstb), .EIYK1nT0oJLxbcxjmodwrC(ds3UaO1QhyfiWT7RZKX23G[0]), .l45qCeMpWMHOXjwYLaHORRE(ds3UaO1QhyfiWT7RZKX23G[1]), .j8SzfGJHmeoXnV9bhAUk40F(ds3UaO1QhyfiWT7RZKX23G[2]), .dMKGmQc7XAB1i3kk2Yk0hH(ds3UaO1QhyfiWT7RZKX23G[3]), .ydI2XfENb2Kl0A3qJMSMBB(tCCvu1nsVn6k0oKnEbNi9E[0]), .nXMdpgmOgBwUAR30aQsd0B(tCCvu1nsVn6k0oKnEbNi9E[1]), .kenMGol9N3qu644VwSIQzD(tCCvu1nsVn6k0oKnEbNi9E[2]), .ovgS7leqdS5z2NH8xqTyeH(tCCvu1nsVn6k0oKnEbNi9E[3]), .eWSF2FqZGP4L33XPl3WfqF(Vc8f45Qo75ucTzy0jKolzE), .KgtpP4p0xLhni3stSN9j2F(ZNDiypKqoG4e82nJIljMu), .bcPgddVda1xlzyptajDlFG(EW7O02E0JPjfI2XYnqHBZB), .kUUVLVsgipRk0xKvCGrGvE(b5ag7OG9oPVwNLOghEh9at) ); assign rQqvnPiwzKpGmREAhe0vF[0] = Vc8f45Qo75ucTzy0jKolzE; assign rQqvnPiwzKpGmREAhe0vF[1] = ZNDiypKqoG4e82nJIljMu; assign rQqvnPiwzKpGmREAhe0vF[2] = EW7O02E0JPjfI2XYnqHBZB; assign rQqvnPiwzKpGmREAhe0vF[3] = b5ag7OG9oPVwNLOghEh9at; assign f2abs_0 = rQqvnPiwzKpGmREAhe0vF[0]; assign f2abs_1 = rQqvnPiwzKpGmREAhe0vF[1]; assign f2abs_2 = rQqvnPiwzKpGmREAhe0vF[2]; assign f2abs_3 = rQqvnPiwzKpGmREAhe0vF[3]; endmodule
