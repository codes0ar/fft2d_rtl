`timescale 1 ns / 1 ns module PxGtD8RdpEuqNR1OqCny8D (v04pHKxyc2sPW047bbyUgE, E7QNJoK4KvAThVFhUlvl2G, l30d1QakAt61ivcMw8sJQE, UKo8akspo4h0jsZ6g712NB, EYQG62ys4E6V8lISAdlW1C, HmVcl5yQin7hEovf3bwNG); parameter integer AddrWidth = 1; parameter integer DataWidth = 1; input v04pHKxyc2sPW047bbyUgE; input signed [DataWidth - 1:0] E7QNJoK4KvAThVFhUlvl2G; input [AddrWidth - 1:0] l30d1QakAt61ivcMw8sJQE; input UKo8akspo4h0jsZ6g712NB; input [AddrWidth - 1:0] EYQG62ys4E6V8lISAdlW1C; output signed [DataWidth - 1:0] HmVcl5yQin7hEovf3bwNG; reg [DataWidth - 1:0] ram [2**AddrWidth - 1:0]; reg [DataWidth - 1:0] data_int; wire QE33642HnVDvOxllaI3KzC; always @(posedge v04pHKxyc2sPW047bbyUgE) begin : PxGtD8RdpEuqNR1OqCny8D_prc if (UKo8akspo4h0jsZ6g712NB == 1'b1) begin ram[l30d1QakAt61ivcMw8sJQE] <= E7QNJoK4KvAThVFhUlvl2G; end data_int <= ram[EYQG62ys4E6V8lISAdlW1C]; end assign HmVcl5yQin7hEovf3bwNG = data_int; endmodule