`timescale 1 ns / 1 ns module UoUhxjuVDf73mwAaAcjVRH (tu9ohhJdK00us7wfvWNQYC, utKZyKAnyhCUOZ6LUagX4D, gA7z08sAKJH0Dq3fae8ZeF, vrNoBb2ZnRj9xKaojUq7EG, b0y2UtjO5W56S6DbL4mEOC, Htw4jhVkz8IRnd9IbKpIUC, y4o9opauBD4PXZzgZLUETHF, yPz5e3igECVkjPPXSkoiHG, z8dRITT2PceChhB9z9EWBC, N7ZKCQ4vfkUB2KkHwgE4GC, PfPBxRXyGunZRp8BSw7dcF, o5kjnQ9W5HT05kz0swOA6QH); input signed [32:0] tu9ohhJdK00us7wfvWNQYC; input signed [32:0] utKZyKAnyhCUOZ6LUagX4D; input signed [32:0] gA7z08sAKJH0Dq3fae8ZeF; input signed [32:0] vrNoBb2ZnRj9xKaojUq7EG; input [17:0] b0y2UtjO5W56S6DbL4mEOC; input [17:0] Htw4jhVkz8IRnd9IbKpIUC; input [17:0] y4o9opauBD4PXZzgZLUETHF; input [17:0] yPz5e3igECVkjPPXSkoiHG; output [17:0] z8dRITT2PceChhB9z9EWBC; output [17:0] N7ZKCQ4vfkUB2KkHwgE4GC; output [17:0] PfPBxRXyGunZRp8BSw7dcF; output [17:0] o5kjnQ9W5HT05kz0swOA6QH; wire [17:0] GHpfOTKsGXKvOOfeyCmWiB [0:3]; wire [17:0] J7L1xgbMCUKJF770vOdvTE; wire [17:0] U4mSpNFxwTaT6m00lo16sD; wire [17:0] PDu13GCvnQyDTshS0WhaTE; wire [17:0] UUaBqOAus1gDnuN8Bmg7wG; wire zx48mBFkrniJrAjwhCL3n; assign GHpfOTKsGXKvOOfeyCmWiB[0] = b0y2UtjO5W56S6DbL4mEOC; assign GHpfOTKsGXKvOOfeyCmWiB[1] = Htw4jhVkz8IRnd9IbKpIUC; assign GHpfOTKsGXKvOOfeyCmWiB[2] = y4o9opauBD4PXZzgZLUETHF; assign GHpfOTKsGXKvOOfeyCmWiB[3] = yPz5e3igECVkjPPXSkoiHG; assign J7L1xgbMCUKJF770vOdvTE = (tu9ohhJdK00us7wfvWNQYC == 33'sh000000000 ? GHpfOTKsGXKvOOfeyCmWiB[0] : (tu9ohhJdK00us7wfvWNQYC == 33'sh000000001 ? GHpfOTKsGXKvOOfeyCmWiB[1] : (tu9ohhJdK00us7wfvWNQYC == 33'sh000000002 ? GHpfOTKsGXKvOOfeyCmWiB[2] : GHpfOTKsGXKvOOfeyCmWiB[3]))); assign z8dRITT2PceChhB9z9EWBC = J7L1xgbMCUKJF770vOdvTE; assign U4mSpNFxwTaT6m00lo16sD = (utKZyKAnyhCUOZ6LUagX4D == 33'sh000000000 ? GHpfOTKsGXKvOOfeyCmWiB[0] : (utKZyKAnyhCUOZ6LUagX4D == 33'sh000000001 ? GHpfOTKsGXKvOOfeyCmWiB[1] : (utKZyKAnyhCUOZ6LUagX4D == 33'sh000000002 ? GHpfOTKsGXKvOOfeyCmWiB[2] : GHpfOTKsGXKvOOfeyCmWiB[3]))); assign N7ZKCQ4vfkUB2KkHwgE4GC = U4mSpNFxwTaT6m00lo16sD; assign PDu13GCvnQyDTshS0WhaTE = (gA7z08sAKJH0Dq3fae8ZeF == 33'sh000000000 ? GHpfOTKsGXKvOOfeyCmWiB[0] : (gA7z08sAKJH0Dq3fae8ZeF == 33'sh000000001 ? GHpfOTKsGXKvOOfeyCmWiB[1] : (gA7z08sAKJH0Dq3fae8ZeF == 33'sh000000002 ? GHpfOTKsGXKvOOfeyCmWiB[2] : GHpfOTKsGXKvOOfeyCmWiB[3]))); assign PfPBxRXyGunZRp8BSw7dcF = PDu13GCvnQyDTshS0WhaTE; assign UUaBqOAus1gDnuN8Bmg7wG = (vrNoBb2ZnRj9xKaojUq7EG == 33'sh000000000 ? GHpfOTKsGXKvOOfeyCmWiB[0] : (vrNoBb2ZnRj9xKaojUq7EG == 33'sh000000001 ? GHpfOTKsGXKvOOfeyCmWiB[1] : (vrNoBb2ZnRj9xKaojUq7EG == 33'sh000000002 ? GHpfOTKsGXKvOOfeyCmWiB[2] : GHpfOTKsGXKvOOfeyCmWiB[3]))); assign o5kjnQ9W5HT05kz0swOA6QH = UUaBqOAus1gDnuN8Bmg7wG; endmodule