`timescale 1 ns / 1 ns module wtU1sSRiRHqGwLWK3NzQmD (v04pHKxyc2sPW047bbyUgE, JAMOfrNHxGSYDF0urqkLN, r3faKvvHpwNbS8m4h6rXSUB, cmM018LKGhcOIt4F15GJS, J5kDQbkAAS4E39jPz9JzwD, PVNB5uj77jMa2DXz4vJtIH, xj2txhdk3kH1ioK0rKOVrG, R6zf5iqRNVEGVBO8egq8kF, mdal5obekPJm0ao7ZiZ4cF, q4mhS1P9mOTwehAXXNmhxF, vyWRmDyKy2RVVIdRBtzV5F, SRoFC9yIIwEIUwYpoyy0QF, wpHiLzmis5ns3l38MddOzE, j963sPBld8mpm71sqcvb8WF, Ic4vfYy6jnxaw8uXI98INH, x2KkW4HKTQgVBmVskDu4RD, g1D8wSsV4Ksuy5G0qxKYMs); input v04pHKxyc2sPW047bbyUgE; input JAMOfrNHxGSYDF0urqkLN; input signed [15:0] r3faKvvHpwNbS8m4h6rXSUB; input signed [15:0] cmM018LKGhcOIt4F15GJS; input signed [15:0] J5kDQbkAAS4E39jPz9JzwD; input signed [15:0] PVNB5uj77jMa2DXz4vJtIH; input xj2txhdk3kH1ioK0rKOVrG; input R6zf5iqRNVEGVBO8egq8kF; output signed [15:0] mdal5obekPJm0ao7ZiZ4cF; output signed [15:0] q4mhS1P9mOTwehAXXNmhxF; output signed [15:0] vyWRmDyKy2RVVIdRBtzV5F; output signed [15:0] SRoFC9yIIwEIUwYpoyy0QF; output signed [15:0] wpHiLzmis5ns3l38MddOzE; output signed [15:0] j963sPBld8mpm71sqcvb8WF; output signed [15:0] Ic4vfYy6jnxaw8uXI98INH; output signed [15:0] x2KkW4HKTQgVBmVskDu4RD; output g1D8wSsV4Ksuy5G0qxKYMs; wire Ebx0yJLDGKevxkqzRPIfvG; wire signed [15:0] YlxyR7WGjsMhhu4Xx4RSSB; reg signed [15:0] XQltXNYzwWy18SM8pDhf8 [0:2]; wire signed [15:0] V1YnWmj1nZzru97DWQqYdE [0:2]; wire signed [15:0] o2uqAyPGPhc9kWis6ko5zF; wire signed [15:0] QGsDAxbcaiCrR87cHhQgZB; reg signed [15:0] TqWcgwsoO3Igmoq6nH36SB [0:2]; wire signed [15:0] pIqvCE2ZCwGFIfCd4j88bF [0:2]; wire signed [15:0] gQqiy8aSxaMx5WfBvElDvC; reg [0:2] c5tyBuJoNrswqnLWL1VV0SB; wire [0:2] mqwYm78twnDBgE5C13tVbH; wire JdpDaA8gpSp0rE35OGZkGE; wire Y7Nx2PyXNCTBUqlHxdhnVC; wire [6:0] u5bboUjXYRZBbt1duYbKTG; wire mir92X5UlUGvLQSXmCuq9; wire hOMBB3qOa4Z6E9dukDYA0F; wire signed [15:0] T5AT5f0lEmroNWkp0Q2apF; wire signed [15:0] y1LfsyMlarAn5fGBZpnPZMF; wire c070CKvbOwMMYffRzNpxjuG; wire pLZcRyd2lMVX3oSoEEblZE; wire [5:0] BZMbpSF4BAilhRWeHczrfC; wire Ax88y9n8GnrKjg0yG0FKzE; wire CosmSfOlF9hl7OPB7KnKvB; wire rFrTP2XEQaUmbjytbnblxB; wire signed [15:0] fLyblCFVFCDbMYyz46VIuE; wire signed [15:0] XaGcqEbv9maW48mW4ZEjUF; wire b93Ikbo3dw8VtPD6KcPt3C; reg signed [15:0] LqbGk6Fit5FCOuam4sOAAD [0:2]; wire signed [15:0] Bi3HF1UTdSkQGHjQ4xRwvF [0:2]; wire signed [15:0] FPJLoZTbR5NUHIeb5WjctB; reg signed [15:0] yLZlCsGdKifpjAYDy4DDED [0:2]; wire signed [15:0] o2lMuceP2Zz2x444DyOgERH [0:2]; wire signed [15:0] j7QbZWviLec2smu8yuKCIPF; reg [0:2] KyQ2PfyWtleyBDhGs5a1gF; wire [0:2] l750CVLudfD6Rvkr3byjjvH; wire pCWATI9lTIGbmXTtLuLAGB; wire signed [15:0] zFuIFDmench8v1O4yXu4jG; wire signed [15:0] dQK1re9uLGxG0WuVGLoXdH; wire kIsHJAwQMWbIiCsXfX1rTG; wire [4:0] yTf5WZbZOLm2uKwJmXk5sG; wire wGlnEfCkRPxniOjCaZH6XG; wire RDvlVEJspE7WkJvNmR8a6C; wire signed [15:0] H8Iagd3fwKKnwcTjUyOkqB; wire signed [15:0] CVOHwOszKLN4rogfAKlMXB; wire DZol1WsbVnSldsei0SiI9E; wire sIaC8spfzCmUwexq8stmB; wire [3:0] zqdZMmoxIs9zmnL4kATVuC; wire a8rK4qdEuNCWHLdYbR2f8; wire O6TgnxqnGk692qEmnZQFTC; wire XfCDnggI1Y1qaMzSOLL0TD; wire signed [15:0] qfBqSs1n7vrUenPHRhvA4E; wire signed [15:0] s1Ni5BKBwo5acvXPnlIkC4D; wire NMWfejbHi1tIjFkylFWDkC; reg signed [15:0] cVMiV2j8qD0P3CVc315hn [0:2]; wire signed [15:0] a9iZ9svlbzlFdVAGUFPTY [0:2]; wire signed [15:0] lyOqtmFbWBeDZLo4tO89VD; reg signed [15:0] u2yic2bBqAL2jFtl9bgNqD [0:2]; wire signed [15:0] rKHf7GW9kd2HwW2mmfwvqC [0:2]; wire signed [15:0] nMEIHp8iZdLbxWoHks1NAB; reg [0:2] qM3kFDhftMVWrl1HT1qB4F; wire [0:2] eHbdLpdf2r0lFYM9BhuRoB; wire v6PtMRDEb2KzMpzXWCSiwkB; wire signed [15:0] HXT3YNFExOHI94Xq9VVUBG; wire signed [15:0] EI1r2DTkmcgS5siR9DUFpG; wire NHkD6RGVcC6B7ibmcHypOC; wire [2:0] u6oVvmCf0f079jLPodlV5B; wire qv4pS1KBm1VYTuOTZHo04F; wire LSv5mOYTPLq5vaIpiVTypC; wire signed [15:0] zsayMT6gR21wpeAixbNYEF; wire signed [15:0] CaTCMDu7mVwW7eYB1tjZ5; wire Ck459KQ1C8vRbine3lrkt; wire DCqZJgzh8RI4wgf1TYRoc; wire [1:0] MCqIdNMOB0Mg1cefHLMjpH; wire j41GwwL8b9NI9l6ZScQ1PbG; wire i8H7HzN3cvjFks6MZ5qaqF; wire SAcShGLK2YZQrWHGqGVvjD; wire signed [15:0] rFr1ZhZNiURIbPFlZaI4kB; wire signed [15:0] gJidztDROiWi1BoJ2KzqKB; wire mm30CTneMiOZJcmmoHkb2D; reg signed [15:0] f69xGE65xXz2LbsT91hgR8G [0:2]; wire signed [15:0] v4gfbuVl5KUcQzK24qqOvB [0:2]; wire signed [15:0] fqWJFy01OVWF8KccC3qB3D; reg signed [15:0] v2G3ZeHqmqPQjfLNmkS0OrG [0:2]; wire signed [15:0] BrQqlwQZdOtmNiJOrBili [0:2]; wire signed [15:0] xQi4zr3ffMHzVne99yIP6E; reg [0:2] k11T3BX1fbEFyiI1W12X7; wire [0:2] VpKk1YVVYHSJ6RsO9pshiB; wire l9QVSAqS6jsMaipvGnosLD; wire signed [15:0] VN3Bh8NuBVl50GFZtWiEND; wire signed [15:0] LEiPXgXUGRZr32PH6jgJWB; wire m0Pt9awzMYrRUb1BRHcMLqG; wire g1oJwDFAtNAcPvLahTlMEB; wire wf5f4XnltnQYt1bEDWEp0F; wire Q7D2KKVRLkwEPktPhyCkSD; wire signed [15:0] LBLHHGcvOnNi88tRjVUMaC; wire signed [15:0] ZKjiEFAXFaCWunBFBNtd0; wire QWAACQosHJOUrDgm1wJeoG; wire hKoHLVfoAgFN4AYEXJutV; wire WgU2KCxd1j6m3EUCPiuf1F; wire y9Hu20tqKGzmg7O1xqeuAZH; wire F9FfK0xrG2zVVJqYJzgfxD; wire xGMN0H1JXsbMHEVz1iuteB; wire signed [15:0] l7IYN7joqiz566PVFOWVRgE; wire signed [15:0] WJrLCpghLrgwyLgXr83JPE; wire NdNevEoWljk83nSbsGDU1C; wire signed [15:0] ZUvkCSPk2wxrRuRb2EYaAH; reg signed [15:0] RAKTymlGVAtDEhqm1mBWKC [0:2]; wire signed [15:0] yyMRtRepkZFuqH6zjb0hbC [0:2]; wire signed [15:0] RclzV3Jlkk5FKKnL0G6JcF; wire signed [15:0] KD169OZrhp2wAmRft0mIM; reg signed [15:0] k9BY0fd7LFxuaZBtnq2NstC [0:2]; wire signed [15:0] mTZgUkGw3710r8TqEV6XWF [0:2]; wire signed [15:0] sueXASR1jeFcZWA77t3pGH; wire signed [15:0] d41CUYvsIlUzO1gIRNNShD; wire signed [15:0] QLKtWBpH0VjEHhv0F6cEGD; wire signed [15:0] LHOKWpKrWmWJXxxXqAj0TH; wire signed [15:0] u9UFtyHKgbvGPJXvb5sSmF; reg signed [15:0] k8gGlV5iKkuIBPqjsMS5KF [0:2]; wire signed [15:0] jVudy6rBy3pL4AAajihjvH [0:2]; wire signed [15:0] DbYwoM2JCYD9mwcRRKmb6G; reg signed [15:0] x9EdsEkQtjpM4w517iGHzC [0:2]; wire signed [15:0] tnuZKwedoQlWAtzBo6aIZB [0:2]; wire signed [15:0] WbySmFpEqdJe6nrpd6KgG; wire signed [15:0] i4y6Td18s9Zr0JbepLQtjC; wire signed [15:0] k3FlrGNoOUOhUgHDIDYGouE; wire signed [15:0] t30W3eeadZl9O9RnQCafyED; wire signed [15:0] flGpcmOyc38fKmqiV5eQvF; wire signed [15:0] CBqrXFTnHQDD2JNQjTxpkH; wire signed [15:0] dYQ3fSOENqw4ZimOQmMMTH; reg signed [15:0] KmuHj4FutgT59Q7oCiggpD [0:2]; wire signed [15:0] UFFCUGMTW5jYs8JEV3j3KC [0:2]; wire signed [15:0] lSTAIQPANZYVi9u1bQJbfC; reg signed [15:0] appAG8sqUT59wY8ObKEssF [0:2]; wire signed [15:0] d21AAbScpxqwLWzuGxj8ajB [0:2]; wire signed [15:0] hh7M8p6TyfjHKgE0YxcN3; wire signed [15:0] FB6nKajjqrTT1538hBpQ9C; wire signed [15:0] XcmpMS0nhYnUzTPGBkEmmF; wire signed [15:0] OAkG388GVoqfAFfrsC3Z3; wire signed [15:0] DP58bSOk4VSBFH6tnqlVTH; wire signed [15:0] oEtRmwXRZkMV2JHZdumYM; wire signed [15:0] ABAJKgUy1j1LH4rwhRtEnG; reg signed [15:0] pISZVQJtPY1M87J4LAx1MB [0:2]; wire signed [15:0] EwyTeOtw0Znxv6WUZIsKtH [0:2]; wire signed [15:0] OTz07QnhICRdmhJUaCsjDD; reg signed [15:0] ufyCKBsm7ZcDMoHa9lVT8B [0:2]; wire signed [15:0] lc0FzXjU6ruJOOuwpT5PQ [0:2]; wire signed [15:0] jnRu1hLACcXOUmEbgPMwFH; wire signed [15:0] NQfJJVPm8CcUv19grKEsZB; wire signed [15:0] k67mERxT6pCrtuCZzqKAJD; wire signed [15:0] lZzpoGgoYZNYjthSDnLuPH; wire signed [15:0] R8WEgTosuCMkRIvxet0i5D; wire signed [15:0] gEaylbF1WXdCOYwXfvD4G; wire signed [15:0] o4iXCc2GyRgQIsHmtR0i8nE; wire signed [15:0] ymBdGOgDsRajoiY9d7TZdC; wire signed [15:0] q8L6STCfvGEzwAAhXRTKviE; wire signed [15:0] EnlAo7K66kKuzHIKWLmc1F; wire signed [15:0] ew3EeLap6s8rXmNrsqaTWH; wire signed [15:0] IPh1M0O3x0ioGlon72MROG; wire signed [15:0] Mt05SNCQbo0cCPNa1yEFyF; wire Z7ZDy0EvwvoCh1zahAqvSF; wire signed [15:0] V7D51SjWfBbpNwnqW3bM8F; reg signed [15:0] f6n0j0rIhtlF1cK7ntOhdG [0:2]; wire signed [15:0] f8PGb7nqRvYgidEKAnbVYCF [0:2]; wire signed [15:0] SvMbkNSHmfXxZeVeRXimM; wire signed [15:0] a9SSaqPU7lUCu5a3eXSIsF; reg signed [15:0] hDe4KgCGLUE2lc3mBRHUGE [0:2]; wire signed [15:0] ZvqDLDMtFPbHpUtzihpbXF [0:2]; wire signed [15:0] qGH0gnrBBGm2QIOAgMsMCH; wire signed [15:0] TyWfuK18qujvo4OtMAdhe; wire signed [15:0] PoiwHvfIvYu5tuiBaljpTF; wire signed [15:0] WdhKnVKybfbzc7shj6T5ID; wire signed [15:0] Z8VgU0v1VN5pqpZolA5AtF; reg signed [15:0] I3TwcvTY4hEZBUKyNKGQYH [0:2]; wire signed [15:0] ltutKZEJ3uAsYBtveZfxN [0:2]; wire signed [15:0] risZnLFYvPBrH1cy6dfHMF; reg signed [15:0] h41dWYc0X3ZAsDk44FMtsTD [0:2]; wire signed [15:0] kZIaatjtNR5S1owTPfmSI [0:2]; wire signed [15:0] y3mUIhc5hpdbI6gB0Klf3MH; wire signed [15:0] UlGc2PVtJa9BNobxUHDxSG; wire signed [15:0] pdTCH0gTlgy9qR74rtvuBE; wire signed [15:0] msLJn85q5aDnigXPSLnA9F; wire signed [15:0] s8tbEDkTdSLkOXc5hVDArH; wire signed [15:0] ACHpp43jQbQJO4HdGlLQ0B; wire signed [15:0] BJNXQzaMpa7r8LYTHlOrBD; reg signed [15:0] UbhppxZFtuRiGSMYxgMT2F [0:2]; wire signed [15:0] rk6XtqxIQmYnoKIvpO9PNH [0:2]; wire signed [15:0] BXAaMHpKzPpYZGFRqoevNE; reg signed [15:0] TGSVeodh4aSh5YMUFsJBpF [0:2]; wire signed [15:0] pKwMCjbBuwX4wlYrJtZeqH [0:2]; wire signed [15:0] czP63K90EaJdtsY9EHZ30D; wire signed [15:0] mxtJaiWQH83FcZ66WqnMiH; wire signed [15:0] MtlWbaE0z2xTCIy368PlWF; wire signed [15:0] Sek0doTmbyRuabtHW5JKgH; wire signed [15:0] h4q2yYljVPy2UhMxEpHXfqG; wire signed [15:0] Ni5CWVNOepdNWeLhPbktyC; wire signed [15:0] oC9IZ8suhbNZiMMpUwYFZE; reg signed [15:0] t1XxIWfdmuGYgMJ14AA5aoF [0:2]; wire signed [15:0] Ed8ZUSDNSkOaxlQSyerJMG [0:2]; wire signed [15:0] lTYYhj3P59f6KeSXhObJAE; reg signed [15:0] u4aeKdZeegD94j2S6reFTD [0:2]; wire signed [15:0] UAnK8iuwkF7gLvWzaOGeMF [0:2]; wire signed [15:0] WawYOEnpsrkHlANz6YaiLG; wire signed [15:0] UwIsRF8C7ejj45D9sxKqgB; wire signed [15:0] XVoYQfnVFtlWlmN3BG5OI; wire signed [15:0] BSsYK6f7nJDXvl3FdklrNE; wire signed [15:0] gGYwPRSrxVg8T85ahN6sK; wire signed [15:0] S6Ue4SxCiz8dBHTO2guOUE; wire signed [15:0] POhLmCr6emegQDte8TzyQ; wire signed [15:0] CyGvS8xQz9obtGAMlB4YwE; reg signed [15:0] G3KM4o4fYtZmkhM463zMWE [0:2]; wire signed [15:0] drYAp2dAOmGqd7jeMIwcRE [0:2]; wire signed [15:0] TAkRd7owTLUvbZtOoRFPtC; wire signed [15:0] imE2eHPyQozGdwpwWRjBLH; reg signed [15:0] RtR9LcVWPsx9vZqDGyBkAB [0:2]; wire signed [15:0] LWmwrv39ujCMpMMcrbgkHC [0:2]; wire signed [15:0] kj4wsLBVI5X3Usybs4WmJH; wire signed [15:0] f3NrgRvCkMfwf1E3PnKtczF; wire signed [15:0] f2XZKbXdctKWPTTQYeLkBWE; wire signed [15:0] f6fgzNt42ufBw7e8PMAUaCB; wire signed [15:0] eYtcM9qmF8eYE3uuCl3HAH; reg signed [15:0] ItzBwvoI4TcHK9g7KBaUVF [0:2]; wire signed [15:0] fk0F6dFxBPneyImhFH4wGG [0:2]; wire signed [15:0] EiKTmNA9gqnqt6QU2ytsGF; reg signed [15:0] VGCjFskQzxD0kIw7klsyNH [0:2]; wire signed [15:0] bsgCRrS7Pvyw5lDPgR03YH [0:2]; wire signed [15:0] i0padod73DFvzROjA4fS2o; wire signed [15:0] mvb8xVo6CcFPFyQu3ctDE; wire signed [15:0] gC05dypmmuscVux3EfDHCD; wire signed [15:0] DxKKPTJNNNGcVbnDyBefdC; wire signed [15:0] z5IVnN9scVD1jMboeUZaZG; wire signed [15:0] y2F62Qir2uvIcDNjqoCgbPG; wire signed [15:0] eJSHu1mAvW9BzbMy0ufWWD; reg signed [15:0] uNvrQvd1Y0KX4XHifVskkH [0:2]; wire signed [15:0] NnZ5dINtMrF9dlFO6TR5yF [0:2]; wire signed [15:0] SNl44VPeKmo2uIh5zCljYE; reg signed [15:0] keFLw9kjnIbUmEw9P3ZHlH [0:2]; wire signed [15:0] TdliLJ6QPHrz19i4ud5ApB [0:2]; wire signed [15:0] AXkTVaeFKW3Cvod76gwXK; wire signed [15:0] PV2GPYF9MTfm6A3VIE3yL; wire signed [15:0] VMMfdu9AIUdQe4XcwZLbSC; wire signed [15:0] BSA6wYLjrd40iGAxWAWPUG; wire signed [15:0] mVsThSJWeEPGLaZQZJ476C; wire signed [15:0] Qjop49qrCNJ2RVI1tmxWK; wire signed [15:0] qtlf3VUxsnDXMsfKMVqqRD; reg signed [15:0] a6YcmlBpfsspWdA41bdAcl [0:2]; wire signed [15:0] LYFiNcEj0dggwMwtkvSMMG [0:2]; wire signed [15:0] g86YyREiAmzs3zk0UOLK0TH; reg signed [15:0] VLlSkvLBi8zwJgPezU50UD [0:2]; wire signed [15:0] VLfdJwrUNkj5uYuSH99PLD [0:2]; wire signed [15:0] KhHmaGBWkoUJ6ybiJ9FvHH; wire signed [15:0] h8QlyPXT2MWg8MvvXSR0uAB; wire signed [15:0] tSs6JTBnsDJvMaRawQm6WF; wire signed [15:0] OJ8T6Dl8xEKAEoVpEfestB; wire signed [15:0] LsWvBUKOjIJIwF6hGU5kRC; wire signed [15:0] E9kfQ0vBTIumIk9ATubhJH; wire signed [15:0] GFkF4uUefeRBOH9Wes3V5D; wire signed [15:0] Tf0EDmJTni9HuTSAYQFT2F; wire signed [15:0] qp9pmnimi6dV0X7tI2Wt6B; wire signed [15:0] Gw5sPQAOzFLVF06eF1AOGF; wire signed [15:0] uO7PvkjtbrbcoMU62rs5JF; wire signed [15:0] qmhLAZZAHFrO09l1zXnPRC; wire signed [15:0] JMtgCMT5TVzyJSn9uILA1; wire signed [15:0] xYJCS7zMCKI1yYR3Bx1XrD; wire signed [15:0] AaqUpSvCGAV1YR86nIsLWH; wire signed [15:0] B58twvtfgVWGK5P29KavtH; wire signed [15:0] qhk6Uhwhppvpssqm7Nh6XE; wire signed [15:0] k3VfrgkD6DWITJL9WW5W4D; wire signed [15:0] pPn6MVGqBLqJ0xzN2WYfFG; wire jNZ4xylBKAANfCL11XNxzB; wire signed [15:0] VWSiqDgxQN9a2J7zRy3p4E; wire signed [15:0] LhqlKpPzANkuN2xC8HYciC; wire signed [15:0] OUMqBzkN19EDa2VTABMa2E; wire signed [15:0] qbEnMIxMUsx8pYkF1gFd7D; wire signed [15:0] A5SQIaNgqW7DcTqQkKRVeD; wire signed [15:0] GaetbCaMty7UkzjqNoYErC; wire signed [15:0] M5AqS9R7rFTkWxwo8io2rH; wire signed [15:0] lcJo4MnEaj41ofRAtLkn4D; wire iyuklaABkAlPLEQPPmVPCD; wire j8MMagsoA5t6IysA2ZD3X4F; wire signed [15:0] aydyoHsGbz0wVGlm34qlsB; wire signed [15:0] H0BpAwmwCivCDsbLQ5qvCC; wire signed [15:0] s1N0USypDrc4xyzxc4XEMr; wire signed [15:0] sZ7bCwrhIAA80IOhzh695; wire dIMToqV6vqVBDOSMMKN0KD; assign Ebx0yJLDGKevxkqzRPIfvG = 1'b0; assign YlxyR7WGjsMhhu4Xx4RSSB = r3faKvvHpwNbS8m4h6rXSUB; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : MczQYJ6MT1pYZD7C1UhQv if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin XQltXNYzwWy18SM8pDhf8[0] <= 16'sb0000000000000000; XQltXNYzwWy18SM8pDhf8[1] <= 16'sb0000000000000000; XQltXNYzwWy18SM8pDhf8[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin XQltXNYzwWy18SM8pDhf8[0] <= 16'sb0000000000000000; XQltXNYzwWy18SM8pDhf8[1] <= 16'sb0000000000000000; XQltXNYzwWy18SM8pDhf8[2] <= 16'sb0000000000000000; end else begin XQltXNYzwWy18SM8pDhf8[0] <= V1YnWmj1nZzru97DWQqYdE[0]; XQltXNYzwWy18SM8pDhf8[1] <= V1YnWmj1nZzru97DWQqYdE[1]; XQltXNYzwWy18SM8pDhf8[2] <= V1YnWmj1nZzru97DWQqYdE[2]; end end end assign o2uqAyPGPhc9kWis6ko5zF = XQltXNYzwWy18SM8pDhf8[2]; assign V1YnWmj1nZzru97DWQqYdE[0] = YlxyR7WGjsMhhu4Xx4RSSB; assign V1YnWmj1nZzru97DWQqYdE[1] = XQltXNYzwWy18SM8pDhf8[0]; assign V1YnWmj1nZzru97DWQqYdE[2] = XQltXNYzwWy18SM8pDhf8[1]; assign QGsDAxbcaiCrR87cHhQgZB = 16'sb0000000000000000; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : xwyxj2YIc64Lxvl4r8S8mG if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin TqWcgwsoO3Igmoq6nH36SB[0] <= 16'sb0000000000000000; TqWcgwsoO3Igmoq6nH36SB[1] <= 16'sb0000000000000000; TqWcgwsoO3Igmoq6nH36SB[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin TqWcgwsoO3Igmoq6nH36SB[0] <= 16'sb0000000000000000; TqWcgwsoO3Igmoq6nH36SB[1] <= 16'sb0000000000000000; TqWcgwsoO3Igmoq6nH36SB[2] <= 16'sb0000000000000000; end else begin TqWcgwsoO3Igmoq6nH36SB[0] <= pIqvCE2ZCwGFIfCd4j88bF[0]; TqWcgwsoO3Igmoq6nH36SB[1] <= pIqvCE2ZCwGFIfCd4j88bF[1]; TqWcgwsoO3Igmoq6nH36SB[2] <= pIqvCE2ZCwGFIfCd4j88bF[2]; end end end assign gQqiy8aSxaMx5WfBvElDvC = TqWcgwsoO3Igmoq6nH36SB[2]; assign pIqvCE2ZCwGFIfCd4j88bF[0] = QGsDAxbcaiCrR87cHhQgZB; assign pIqvCE2ZCwGFIfCd4j88bF[1] = TqWcgwsoO3Igmoq6nH36SB[0]; assign pIqvCE2ZCwGFIfCd4j88bF[2] = TqWcgwsoO3Igmoq6nH36SB[1]; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : L1HBH8O5DRbGBa9XvBX70C if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin c5tyBuJoNrswqnLWL1VV0SB[0] <= 1'b0; c5tyBuJoNrswqnLWL1VV0SB[1] <= 1'b0; c5tyBuJoNrswqnLWL1VV0SB[2] <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin c5tyBuJoNrswqnLWL1VV0SB[0] <= 1'b0; c5tyBuJoNrswqnLWL1VV0SB[1] <= 1'b0; c5tyBuJoNrswqnLWL1VV0SB[2] <= 1'b0; end else begin c5tyBuJoNrswqnLWL1VV0SB[0] <= mqwYm78twnDBgE5C13tVbH[0]; c5tyBuJoNrswqnLWL1VV0SB[1] <= mqwYm78twnDBgE5C13tVbH[1]; c5tyBuJoNrswqnLWL1VV0SB[2] <= mqwYm78twnDBgE5C13tVbH[2]; end end end assign JdpDaA8gpSp0rE35OGZkGE = c5tyBuJoNrswqnLWL1VV0SB[2]; assign mqwYm78twnDBgE5C13tVbH[0] = xj2txhdk3kH1ioK0rKOVrG; assign mqwYm78twnDBgE5C13tVbH[1] = c5tyBuJoNrswqnLWL1VV0SB[0]; assign mqwYm78twnDBgE5C13tVbH[2] = c5tyBuJoNrswqnLWL1VV0SB[1]; Jwp87To0uCqWGVPIwhN8ED RGbrDjFygXYGvFvOLlE8vD (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .Y7Nx2PyXNCTBUqlHxdhnVC(Y7Nx2PyXNCTBUqlHxdhnVC), .w9tDlZkclLF2jmOsqVKqWE(Y7Nx2PyXNCTBUqlHxdhnVC), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .u5bboUjXYRZBbt1duYbKTG(u5bboUjXYRZBbt1duYbKTG), .mir92X5UlUGvLQSXmCuq9(mir92X5UlUGvLQSXmCuq9), .hOMBB3qOa4Z6E9dukDYA0F(hOMBB3qOa4Z6E9dukDYA0F) ); YBvtcUvICoqzwziatY4vk U3WFM5mS8kDgJTOIhMNlWE (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .o2uqAyPGPhc9kWis6ko5zF(o2uqAyPGPhc9kWis6ko5zF), .gQqiy8aSxaMx5WfBvElDvC(gQqiy8aSxaMx5WfBvElDvC), .JdpDaA8gpSp0rE35OGZkGE(JdpDaA8gpSp0rE35OGZkGE), .u5bboUjXYRZBbt1duYbKTG(u5bboUjXYRZBbt1duYbKTG), .mir92X5UlUGvLQSXmCuq9(mir92X5UlUGvLQSXmCuq9), .hOMBB3qOa4Z6E9dukDYA0F(hOMBB3qOa4Z6E9dukDYA0F), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .T5AT5f0lEmroNWkp0Q2apF(T5AT5f0lEmroNWkp0Q2apF), .y1LfsyMlarAn5fGBZpnPZMF(y1LfsyMlarAn5fGBZpnPZMF), .c070CKvbOwMMYffRzNpxjuG(c070CKvbOwMMYffRzNpxjuG), .Y7Nx2PyXNCTBUqlHxdhnVC(Y7Nx2PyXNCTBUqlHxdhnVC) ); e61uBMMOD8obk5m2QBgMSL IluUflSX1mHXxHZ5bHGXV (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .c070CKvbOwMMYffRzNpxjuG(c070CKvbOwMMYffRzNpxjuG), .pLZcRyd2lMVX3oSoEEblZE(pLZcRyd2lMVX3oSoEEblZE), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .BZMbpSF4BAilhRWeHczrfC(BZMbpSF4BAilhRWeHczrfC), .Ax88y9n8GnrKjg0yG0FKzE(Ax88y9n8GnrKjg0yG0FKzE), .CosmSfOlF9hl7OPB7KnKvB(CosmSfOlF9hl7OPB7KnKvB), .rFrTP2XEQaUmbjytbnblxB(rFrTP2XEQaUmbjytbnblxB) ); w8xdha0uhSMB2MNkwcBaRdB eDGyALcRao2ynBOyHNXQBC (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .T5AT5f0lEmroNWkp0Q2apF(T5AT5f0lEmroNWkp0Q2apF), .y1LfsyMlarAn5fGBZpnPZMF(y1LfsyMlarAn5fGBZpnPZMF), .c070CKvbOwMMYffRzNpxjuG(c070CKvbOwMMYffRzNpxjuG), .BZMbpSF4BAilhRWeHczrfC(BZMbpSF4BAilhRWeHczrfC), .Ax88y9n8GnrKjg0yG0FKzE(Ax88y9n8GnrKjg0yG0FKzE), .CosmSfOlF9hl7OPB7KnKvB(CosmSfOlF9hl7OPB7KnKvB), .rFrTP2XEQaUmbjytbnblxB(rFrTP2XEQaUmbjytbnblxB), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .fLyblCFVFCDbMYyz46VIuE(fLyblCFVFCDbMYyz46VIuE), .XaGcqEbv9maW48mW4ZEjUF(XaGcqEbv9maW48mW4ZEjUF), .b93Ikbo3dw8VtPD6KcPt3C(b93Ikbo3dw8VtPD6KcPt3C), .pLZcRyd2lMVX3oSoEEblZE(pLZcRyd2lMVX3oSoEEblZE) ); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : s2CWr6rrksK4W7N0omU97HD if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin LqbGk6Fit5FCOuam4sOAAD[0] <= 16'sb0000000000000000; LqbGk6Fit5FCOuam4sOAAD[1] <= 16'sb0000000000000000; LqbGk6Fit5FCOuam4sOAAD[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin LqbGk6Fit5FCOuam4sOAAD[0] <= 16'sb0000000000000000; LqbGk6Fit5FCOuam4sOAAD[1] <= 16'sb0000000000000000; LqbGk6Fit5FCOuam4sOAAD[2] <= 16'sb0000000000000000; end else begin LqbGk6Fit5FCOuam4sOAAD[0] <= Bi3HF1UTdSkQGHjQ4xRwvF[0]; LqbGk6Fit5FCOuam4sOAAD[1] <= Bi3HF1UTdSkQGHjQ4xRwvF[1]; LqbGk6Fit5FCOuam4sOAAD[2] <= Bi3HF1UTdSkQGHjQ4xRwvF[2]; end end end assign FPJLoZTbR5NUHIeb5WjctB = LqbGk6Fit5FCOuam4sOAAD[2]; assign Bi3HF1UTdSkQGHjQ4xRwvF[0] = fLyblCFVFCDbMYyz46VIuE; assign Bi3HF1UTdSkQGHjQ4xRwvF[1] = LqbGk6Fit5FCOuam4sOAAD[0]; assign Bi3HF1UTdSkQGHjQ4xRwvF[2] = LqbGk6Fit5FCOuam4sOAAD[1]; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : k1Zsi6BUVrSUjLbIYwh26G if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin yLZlCsGdKifpjAYDy4DDED[0] <= 16'sb0000000000000000; yLZlCsGdKifpjAYDy4DDED[1] <= 16'sb0000000000000000; yLZlCsGdKifpjAYDy4DDED[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin yLZlCsGdKifpjAYDy4DDED[0] <= 16'sb0000000000000000; yLZlCsGdKifpjAYDy4DDED[1] <= 16'sb0000000000000000; yLZlCsGdKifpjAYDy4DDED[2] <= 16'sb0000000000000000; end else begin yLZlCsGdKifpjAYDy4DDED[0] <= o2lMuceP2Zz2x444DyOgERH[0]; yLZlCsGdKifpjAYDy4DDED[1] <= o2lMuceP2Zz2x444DyOgERH[1]; yLZlCsGdKifpjAYDy4DDED[2] <= o2lMuceP2Zz2x444DyOgERH[2]; end end end assign j7QbZWviLec2smu8yuKCIPF = yLZlCsGdKifpjAYDy4DDED[2]; assign o2lMuceP2Zz2x444DyOgERH[0] = XaGcqEbv9maW48mW4ZEjUF; assign o2lMuceP2Zz2x444DyOgERH[1] = yLZlCsGdKifpjAYDy4DDED[0]; assign o2lMuceP2Zz2x444DyOgERH[2] = yLZlCsGdKifpjAYDy4DDED[1]; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : TPi3Fu9uFLztbkFwa0H53D if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin KyQ2PfyWtleyBDhGs5a1gF[0] <= 1'b0; KyQ2PfyWtleyBDhGs5a1gF[1] <= 1'b0; KyQ2PfyWtleyBDhGs5a1gF[2] <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin KyQ2PfyWtleyBDhGs5a1gF[0] <= 1'b0; KyQ2PfyWtleyBDhGs5a1gF[1] <= 1'b0; KyQ2PfyWtleyBDhGs5a1gF[2] <= 1'b0; end else begin KyQ2PfyWtleyBDhGs5a1gF[0] <= l750CVLudfD6Rvkr3byjjvH[0]; KyQ2PfyWtleyBDhGs5a1gF[1] <= l750CVLudfD6Rvkr3byjjvH[1]; KyQ2PfyWtleyBDhGs5a1gF[2] <= l750CVLudfD6Rvkr3byjjvH[2]; end end end assign pCWATI9lTIGbmXTtLuLAGB = KyQ2PfyWtleyBDhGs5a1gF[2]; assign l750CVLudfD6Rvkr3byjjvH[0] = b93Ikbo3dw8VtPD6KcPt3C; assign l750CVLudfD6Rvkr3byjjvH[1] = KyQ2PfyWtleyBDhGs5a1gF[0]; assign l750CVLudfD6Rvkr3byjjvH[2] = KyQ2PfyWtleyBDhGs5a1gF[1]; DxhqsB4bELEu0qDWWrg1F qTfyhdbQzAKcKbDpRJj8yG (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .b93Ikbo3dw8VtPD6KcPt3C(b93Ikbo3dw8VtPD6KcPt3C), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .zFuIFDmench8v1O4yXu4jG(zFuIFDmench8v1O4yXu4jG), .dQK1re9uLGxG0WuVGLoXdH(dQK1re9uLGxG0WuVGLoXdH) ); CF4YZpD8T3bZDeoOS74nFB JSNmXQ0YI7nAzGfsGLG1UC (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .kIsHJAwQMWbIiCsXfX1rTG(kIsHJAwQMWbIiCsXfX1rTG), .DKGIysOp4cb2Wy4ifYHB8D(kIsHJAwQMWbIiCsXfX1rTG), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .yTf5WZbZOLm2uKwJmXk5sG(yTf5WZbZOLm2uKwJmXk5sG), .wGlnEfCkRPxniOjCaZH6XG(wGlnEfCkRPxniOjCaZH6XG), .RDvlVEJspE7WkJvNmR8a6C(RDvlVEJspE7WkJvNmR8a6C) ); dhkIZRHmRjY0Gsp76QLRYH rKXyl8hgTMym1rEDLsJaOB (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .FPJLoZTbR5NUHIeb5WjctB(FPJLoZTbR5NUHIeb5WjctB), .j7QbZWviLec2smu8yuKCIPF(j7QbZWviLec2smu8yuKCIPF), .pCWATI9lTIGbmXTtLuLAGB(pCWATI9lTIGbmXTtLuLAGB), .yTf5WZbZOLm2uKwJmXk5sG(yTf5WZbZOLm2uKwJmXk5sG), .wGlnEfCkRPxniOjCaZH6XG(wGlnEfCkRPxniOjCaZH6XG), .zFuIFDmench8v1O4yXu4jG(zFuIFDmench8v1O4yXu4jG), .dQK1re9uLGxG0WuVGLoXdH(dQK1re9uLGxG0WuVGLoXdH), .RDvlVEJspE7WkJvNmR8a6C(RDvlVEJspE7WkJvNmR8a6C), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .H8Iagd3fwKKnwcTjUyOkqB(H8Iagd3fwKKnwcTjUyOkqB), .CVOHwOszKLN4rogfAKlMXB(CVOHwOszKLN4rogfAKlMXB), .DZol1WsbVnSldsei0SiI9E(DZol1WsbVnSldsei0SiI9E), .kIsHJAwQMWbIiCsXfX1rTG(kIsHJAwQMWbIiCsXfX1rTG) ); T1MCYG31QHzAKthZjSBalB z962IOrouyDUWLniu10oD3C (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .DZol1WsbVnSldsei0SiI9E(DZol1WsbVnSldsei0SiI9E), .sIaC8spfzCmUwexq8stmB(sIaC8spfzCmUwexq8stmB), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .zqdZMmoxIs9zmnL4kATVuC(zqdZMmoxIs9zmnL4kATVuC), .a8rK4qdEuNCWHLdYbR2f8(a8rK4qdEuNCWHLdYbR2f8), .O6TgnxqnGk692qEmnZQFTC(O6TgnxqnGk692qEmnZQFTC), .XfCDnggI1Y1qaMzSOLL0TD(XfCDnggI1Y1qaMzSOLL0TD) ); m3456FzWsQW24e0Gmggh3HD onkga9gnAWHYkWnfgU4ydB (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .H8Iagd3fwKKnwcTjUyOkqB(H8Iagd3fwKKnwcTjUyOkqB), .CVOHwOszKLN4rogfAKlMXB(CVOHwOszKLN4rogfAKlMXB), .DZol1WsbVnSldsei0SiI9E(DZol1WsbVnSldsei0SiI9E), .zqdZMmoxIs9zmnL4kATVuC(zqdZMmoxIs9zmnL4kATVuC), .a8rK4qdEuNCWHLdYbR2f8(a8rK4qdEuNCWHLdYbR2f8), .O6TgnxqnGk692qEmnZQFTC(O6TgnxqnGk692qEmnZQFTC), .XfCDnggI1Y1qaMzSOLL0TD(XfCDnggI1Y1qaMzSOLL0TD), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .qfBqSs1n7vrUenPHRhvA4E(qfBqSs1n7vrUenPHRhvA4E), .s1Ni5BKBwo5acvXPnlIkC4D(s1Ni5BKBwo5acvXPnlIkC4D), .NMWfejbHi1tIjFkylFWDkC(NMWfejbHi1tIjFkylFWDkC), .sIaC8spfzCmUwexq8stmB(sIaC8spfzCmUwexq8stmB) ); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : IBmSJmjQmOQZECy1AykU1D if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin cVMiV2j8qD0P3CVc315hn[0] <= 16'sb0000000000000000; cVMiV2j8qD0P3CVc315hn[1] <= 16'sb0000000000000000; cVMiV2j8qD0P3CVc315hn[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin cVMiV2j8qD0P3CVc315hn[0] <= 16'sb0000000000000000; cVMiV2j8qD0P3CVc315hn[1] <= 16'sb0000000000000000; cVMiV2j8qD0P3CVc315hn[2] <= 16'sb0000000000000000; end else begin cVMiV2j8qD0P3CVc315hn[0] <= a9iZ9svlbzlFdVAGUFPTY[0]; cVMiV2j8qD0P3CVc315hn[1] <= a9iZ9svlbzlFdVAGUFPTY[1]; cVMiV2j8qD0P3CVc315hn[2] <= a9iZ9svlbzlFdVAGUFPTY[2]; end end end assign lyOqtmFbWBeDZLo4tO89VD = cVMiV2j8qD0P3CVc315hn[2]; assign a9iZ9svlbzlFdVAGUFPTY[0] = qfBqSs1n7vrUenPHRhvA4E; assign a9iZ9svlbzlFdVAGUFPTY[1] = cVMiV2j8qD0P3CVc315hn[0]; assign a9iZ9svlbzlFdVAGUFPTY[2] = cVMiV2j8qD0P3CVc315hn[1]; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : VNPcEW4KZxpAtEz0DCT8vD if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin u2yic2bBqAL2jFtl9bgNqD[0] <= 16'sb0000000000000000; u2yic2bBqAL2jFtl9bgNqD[1] <= 16'sb0000000000000000; u2yic2bBqAL2jFtl9bgNqD[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin u2yic2bBqAL2jFtl9bgNqD[0] <= 16'sb0000000000000000; u2yic2bBqAL2jFtl9bgNqD[1] <= 16'sb0000000000000000; u2yic2bBqAL2jFtl9bgNqD[2] <= 16'sb0000000000000000; end else begin u2yic2bBqAL2jFtl9bgNqD[0] <= rKHf7GW9kd2HwW2mmfwvqC[0]; u2yic2bBqAL2jFtl9bgNqD[1] <= rKHf7GW9kd2HwW2mmfwvqC[1]; u2yic2bBqAL2jFtl9bgNqD[2] <= rKHf7GW9kd2HwW2mmfwvqC[2]; end end end assign nMEIHp8iZdLbxWoHks1NAB = u2yic2bBqAL2jFtl9bgNqD[2]; assign rKHf7GW9kd2HwW2mmfwvqC[0] = s1Ni5BKBwo5acvXPnlIkC4D; assign rKHf7GW9kd2HwW2mmfwvqC[1] = u2yic2bBqAL2jFtl9bgNqD[0]; assign rKHf7GW9kd2HwW2mmfwvqC[2] = u2yic2bBqAL2jFtl9bgNqD[1]; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : t8uWAeIAh3IMbN9UNxoYBKD if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin qM3kFDhftMVWrl1HT1qB4F[0] <= 1'b0; qM3kFDhftMVWrl1HT1qB4F[1] <= 1'b0; qM3kFDhftMVWrl1HT1qB4F[2] <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin qM3kFDhftMVWrl1HT1qB4F[0] <= 1'b0; qM3kFDhftMVWrl1HT1qB4F[1] <= 1'b0; qM3kFDhftMVWrl1HT1qB4F[2] <= 1'b0; end else begin qM3kFDhftMVWrl1HT1qB4F[0] <= eHbdLpdf2r0lFYM9BhuRoB[0]; qM3kFDhftMVWrl1HT1qB4F[1] <= eHbdLpdf2r0lFYM9BhuRoB[1]; qM3kFDhftMVWrl1HT1qB4F[2] <= eHbdLpdf2r0lFYM9BhuRoB[2]; end end end assign v6PtMRDEb2KzMpzXWCSiwkB = qM3kFDhftMVWrl1HT1qB4F[2]; assign eHbdLpdf2r0lFYM9BhuRoB[0] = NMWfejbHi1tIjFkylFWDkC; assign eHbdLpdf2r0lFYM9BhuRoB[1] = qM3kFDhftMVWrl1HT1qB4F[0]; assign eHbdLpdf2r0lFYM9BhuRoB[2] = qM3kFDhftMVWrl1HT1qB4F[1]; YWcbaK4GTT05DhR2SHpPIG mYbRzIp6fh5UU50NIPMlqE (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .NMWfejbHi1tIjFkylFWDkC(NMWfejbHi1tIjFkylFWDkC), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .HXT3YNFExOHI94Xq9VVUBG(HXT3YNFExOHI94Xq9VVUBG), .EI1r2DTkmcgS5siR9DUFpG(EI1r2DTkmcgS5siR9DUFpG) ); wxj68aRjPtPccZFhxDpbaE K59tEegFJMrdmJIuWBI7q (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .NHkD6RGVcC6B7ibmcHypOC(NHkD6RGVcC6B7ibmcHypOC), .n6CG7K4rgMGw86VJoKnfuOD(NHkD6RGVcC6B7ibmcHypOC), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .u6oVvmCf0f079jLPodlV5B(u6oVvmCf0f079jLPodlV5B), .qv4pS1KBm1VYTuOTZHo04F(qv4pS1KBm1VYTuOTZHo04F), .LSv5mOYTPLq5vaIpiVTypC(LSv5mOYTPLq5vaIpiVTypC) ); nZi1Oyqdh8BgpskwTUd8GE YGfiJxj5wy9c9fxm8qBmQC (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .lyOqtmFbWBeDZLo4tO89VD(lyOqtmFbWBeDZLo4tO89VD), .nMEIHp8iZdLbxWoHks1NAB(nMEIHp8iZdLbxWoHks1NAB), .v6PtMRDEb2KzMpzXWCSiwkB(v6PtMRDEb2KzMpzXWCSiwkB), .u6oVvmCf0f079jLPodlV5B(u6oVvmCf0f079jLPodlV5B), .qv4pS1KBm1VYTuOTZHo04F(qv4pS1KBm1VYTuOTZHo04F), .HXT3YNFExOHI94Xq9VVUBG(HXT3YNFExOHI94Xq9VVUBG), .EI1r2DTkmcgS5siR9DUFpG(EI1r2DTkmcgS5siR9DUFpG), .LSv5mOYTPLq5vaIpiVTypC(LSv5mOYTPLq5vaIpiVTypC), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .zsayMT6gR21wpeAixbNYEF(zsayMT6gR21wpeAixbNYEF), .CaTCMDu7mVwW7eYB1tjZ5(CaTCMDu7mVwW7eYB1tjZ5), .Ck459KQ1C8vRbine3lrkt(Ck459KQ1C8vRbine3lrkt), .NHkD6RGVcC6B7ibmcHypOC(NHkD6RGVcC6B7ibmcHypOC) ); J2jBxTkCbwexjojaErwtkC BoxmA9gUrcoGKTr1WWdljB (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .Ck459KQ1C8vRbine3lrkt(Ck459KQ1C8vRbine3lrkt), .DCqZJgzh8RI4wgf1TYRoc(DCqZJgzh8RI4wgf1TYRoc), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .MCqIdNMOB0Mg1cefHLMjpH(MCqIdNMOB0Mg1cefHLMjpH), .j41GwwL8b9NI9l6ZScQ1PbG(j41GwwL8b9NI9l6ZScQ1PbG), .i8H7HzN3cvjFks6MZ5qaqF(i8H7HzN3cvjFks6MZ5qaqF), .SAcShGLK2YZQrWHGqGVvjD(SAcShGLK2YZQrWHGqGVvjD) ); Pe7UEMNFrda6tk7SdC5JqB v4tQ5NbkvrLEoEVGS2hwT8F (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .zsayMT6gR21wpeAixbNYEF(zsayMT6gR21wpeAixbNYEF), .CaTCMDu7mVwW7eYB1tjZ5(CaTCMDu7mVwW7eYB1tjZ5), .Ck459KQ1C8vRbine3lrkt(Ck459KQ1C8vRbine3lrkt), .MCqIdNMOB0Mg1cefHLMjpH(MCqIdNMOB0Mg1cefHLMjpH), .j41GwwL8b9NI9l6ZScQ1PbG(j41GwwL8b9NI9l6ZScQ1PbG), .i8H7HzN3cvjFks6MZ5qaqF(i8H7HzN3cvjFks6MZ5qaqF), .SAcShGLK2YZQrWHGqGVvjD(SAcShGLK2YZQrWHGqGVvjD), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .rFr1ZhZNiURIbPFlZaI4kB(rFr1ZhZNiURIbPFlZaI4kB), .gJidztDROiWi1BoJ2KzqKB(gJidztDROiWi1BoJ2KzqKB), .mm30CTneMiOZJcmmoHkb2D(mm30CTneMiOZJcmmoHkb2D), .DCqZJgzh8RI4wgf1TYRoc(DCqZJgzh8RI4wgf1TYRoc) ); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : QtzxgwI206U33aXvIkKdwD if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin f69xGE65xXz2LbsT91hgR8G[0] <= 16'sb0000000000000000; f69xGE65xXz2LbsT91hgR8G[1] <= 16'sb0000000000000000; f69xGE65xXz2LbsT91hgR8G[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin f69xGE65xXz2LbsT91hgR8G[0] <= 16'sb0000000000000000; f69xGE65xXz2LbsT91hgR8G[1] <= 16'sb0000000000000000; f69xGE65xXz2LbsT91hgR8G[2] <= 16'sb0000000000000000; end else begin f69xGE65xXz2LbsT91hgR8G[0] <= v4gfbuVl5KUcQzK24qqOvB[0]; f69xGE65xXz2LbsT91hgR8G[1] <= v4gfbuVl5KUcQzK24qqOvB[1]; f69xGE65xXz2LbsT91hgR8G[2] <= v4gfbuVl5KUcQzK24qqOvB[2]; end end end assign fqWJFy01OVWF8KccC3qB3D = f69xGE65xXz2LbsT91hgR8G[2]; assign v4gfbuVl5KUcQzK24qqOvB[0] = rFr1ZhZNiURIbPFlZaI4kB; assign v4gfbuVl5KUcQzK24qqOvB[1] = f69xGE65xXz2LbsT91hgR8G[0]; assign v4gfbuVl5KUcQzK24qqOvB[2] = f69xGE65xXz2LbsT91hgR8G[1]; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : awX33YTQEl2OxkV2HHm04D if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin v2G3ZeHqmqPQjfLNmkS0OrG[0] <= 16'sb0000000000000000; v2G3ZeHqmqPQjfLNmkS0OrG[1] <= 16'sb0000000000000000; v2G3ZeHqmqPQjfLNmkS0OrG[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin v2G3ZeHqmqPQjfLNmkS0OrG[0] <= 16'sb0000000000000000; v2G3ZeHqmqPQjfLNmkS0OrG[1] <= 16'sb0000000000000000; v2G3ZeHqmqPQjfLNmkS0OrG[2] <= 16'sb0000000000000000; end else begin v2G3ZeHqmqPQjfLNmkS0OrG[0] <= BrQqlwQZdOtmNiJOrBili[0]; v2G3ZeHqmqPQjfLNmkS0OrG[1] <= BrQqlwQZdOtmNiJOrBili[1]; v2G3ZeHqmqPQjfLNmkS0OrG[2] <= BrQqlwQZdOtmNiJOrBili[2]; end end end assign xQi4zr3ffMHzVne99yIP6E = v2G3ZeHqmqPQjfLNmkS0OrG[2]; assign BrQqlwQZdOtmNiJOrBili[0] = gJidztDROiWi1BoJ2KzqKB; assign BrQqlwQZdOtmNiJOrBili[1] = v2G3ZeHqmqPQjfLNmkS0OrG[0]; assign BrQqlwQZdOtmNiJOrBili[2] = v2G3ZeHqmqPQjfLNmkS0OrG[1]; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : wroVmvZXsLz1H55Ur0PrpB if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin k11T3BX1fbEFyiI1W12X7[0] <= 1'b0; k11T3BX1fbEFyiI1W12X7[1] <= 1'b0; k11T3BX1fbEFyiI1W12X7[2] <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin k11T3BX1fbEFyiI1W12X7[0] <= 1'b0; k11T3BX1fbEFyiI1W12X7[1] <= 1'b0; k11T3BX1fbEFyiI1W12X7[2] <= 1'b0; end else begin k11T3BX1fbEFyiI1W12X7[0] <= VpKk1YVVYHSJ6RsO9pshiB[0]; k11T3BX1fbEFyiI1W12X7[1] <= VpKk1YVVYHSJ6RsO9pshiB[1]; k11T3BX1fbEFyiI1W12X7[2] <= VpKk1YVVYHSJ6RsO9pshiB[2]; end end end assign l9QVSAqS6jsMaipvGnosLD = k11T3BX1fbEFyiI1W12X7[2]; assign VpKk1YVVYHSJ6RsO9pshiB[0] = mm30CTneMiOZJcmmoHkb2D; assign VpKk1YVVYHSJ6RsO9pshiB[1] = k11T3BX1fbEFyiI1W12X7[0]; assign VpKk1YVVYHSJ6RsO9pshiB[2] = k11T3BX1fbEFyiI1W12X7[1]; pfUwRLxGLn8DQv6jMCaY3E MwRmE5s9T5vHnHIPrZpBXG (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .mm30CTneMiOZJcmmoHkb2D(mm30CTneMiOZJcmmoHkb2D), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .VN3Bh8NuBVl50GFZtWiEND(VN3Bh8NuBVl50GFZtWiEND), .LEiPXgXUGRZr32PH6jgJWB(LEiPXgXUGRZr32PH6jgJWB) ); CQ8VhzX2aZDdqpzcRKBClF g76zMlLb1BXfd6xhVWKwvIF (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .m0Pt9awzMYrRUb1BRHcMLqG(m0Pt9awzMYrRUb1BRHcMLqG), .o3XsAkfAYoavjVukPhwjwlC(m0Pt9awzMYrRUb1BRHcMLqG), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .g1oJwDFAtNAcPvLahTlMEB(g1oJwDFAtNAcPvLahTlMEB), .wf5f4XnltnQYt1bEDWEp0F(wf5f4XnltnQYt1bEDWEp0F), .Q7D2KKVRLkwEPktPhyCkSD(Q7D2KKVRLkwEPktPhyCkSD) ); RQbqWmk4vKJGwrZzxhzMXF lHIW1e1kbWo3lWzndJPvuB (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .fqWJFy01OVWF8KccC3qB3D(fqWJFy01OVWF8KccC3qB3D), .xQi4zr3ffMHzVne99yIP6E(xQi4zr3ffMHzVne99yIP6E), .l9QVSAqS6jsMaipvGnosLD(l9QVSAqS6jsMaipvGnosLD), .g1oJwDFAtNAcPvLahTlMEB(g1oJwDFAtNAcPvLahTlMEB), .wf5f4XnltnQYt1bEDWEp0F(wf5f4XnltnQYt1bEDWEp0F), .VN3Bh8NuBVl50GFZtWiEND(VN3Bh8NuBVl50GFZtWiEND), .LEiPXgXUGRZr32PH6jgJWB(LEiPXgXUGRZr32PH6jgJWB), .Q7D2KKVRLkwEPktPhyCkSD(Q7D2KKVRLkwEPktPhyCkSD), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .LBLHHGcvOnNi88tRjVUMaC(LBLHHGcvOnNi88tRjVUMaC), .ZKjiEFAXFaCWunBFBNtd0(ZKjiEFAXFaCWunBFBNtd0), .QWAACQosHJOUrDgm1wJeoG(QWAACQosHJOUrDgm1wJeoG), .m0Pt9awzMYrRUb1BRHcMLqG(m0Pt9awzMYrRUb1BRHcMLqG) ); rUdEDJxz9hCFSCEPZfs0dH JJ0nVDqYyN2uYKveWElyMB (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .QWAACQosHJOUrDgm1wJeoG(QWAACQosHJOUrDgm1wJeoG), .hKoHLVfoAgFN4AYEXJutV(hKoHLVfoAgFN4AYEXJutV), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .WgU2KCxd1j6m3EUCPiuf1F(WgU2KCxd1j6m3EUCPiuf1F), .y9Hu20tqKGzmg7O1xqeuAZH(y9Hu20tqKGzmg7O1xqeuAZH), .F9FfK0xrG2zVVJqYJzgfxD(F9FfK0xrG2zVVJqYJzgfxD), .xGMN0H1JXsbMHEVz1iuteB(xGMN0H1JXsbMHEVz1iuteB) ); eCat9Y3EIg6dfvYxFCPRtH xq2LeFrsREQ5RUVqGKULHE (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .LBLHHGcvOnNi88tRjVUMaC(LBLHHGcvOnNi88tRjVUMaC), .ZKjiEFAXFaCWunBFBNtd0(ZKjiEFAXFaCWunBFBNtd0), .QWAACQosHJOUrDgm1wJeoG(QWAACQosHJOUrDgm1wJeoG), .WgU2KCxd1j6m3EUCPiuf1F(WgU2KCxd1j6m3EUCPiuf1F), .y9Hu20tqKGzmg7O1xqeuAZH(y9Hu20tqKGzmg7O1xqeuAZH), .F9FfK0xrG2zVVJqYJzgfxD(F9FfK0xrG2zVVJqYJzgfxD), .xGMN0H1JXsbMHEVz1iuteB(xGMN0H1JXsbMHEVz1iuteB), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .l7IYN7joqiz566PVFOWVRgE(l7IYN7joqiz566PVFOWVRgE), .WJrLCpghLrgwyLgXr83JPE(WJrLCpghLrgwyLgXr83JPE), .NdNevEoWljk83nSbsGDU1C(NdNevEoWljk83nSbsGDU1C), .hKoHLVfoAgFN4AYEXJutV(hKoHLVfoAgFN4AYEXJutV) ); assign ZUvkCSPk2wxrRuRb2EYaAH = cmM018LKGhcOIt4F15GJS; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : z8NMcVNSFzdoHNpSsC5DBLF if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin RAKTymlGVAtDEhqm1mBWKC[0] <= 16'sb0000000000000000; RAKTymlGVAtDEhqm1mBWKC[1] <= 16'sb0000000000000000; RAKTymlGVAtDEhqm1mBWKC[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin RAKTymlGVAtDEhqm1mBWKC[0] <= 16'sb0000000000000000; RAKTymlGVAtDEhqm1mBWKC[1] <= 16'sb0000000000000000; RAKTymlGVAtDEhqm1mBWKC[2] <= 16'sb0000000000000000; end else begin RAKTymlGVAtDEhqm1mBWKC[0] <= yyMRtRepkZFuqH6zjb0hbC[0]; RAKTymlGVAtDEhqm1mBWKC[1] <= yyMRtRepkZFuqH6zjb0hbC[1]; RAKTymlGVAtDEhqm1mBWKC[2] <= yyMRtRepkZFuqH6zjb0hbC[2]; end end end assign RclzV3Jlkk5FKKnL0G6JcF = RAKTymlGVAtDEhqm1mBWKC[2]; assign yyMRtRepkZFuqH6zjb0hbC[0] = ZUvkCSPk2wxrRuRb2EYaAH; assign yyMRtRepkZFuqH6zjb0hbC[1] = RAKTymlGVAtDEhqm1mBWKC[0]; assign yyMRtRepkZFuqH6zjb0hbC[2] = RAKTymlGVAtDEhqm1mBWKC[1]; assign KD169OZrhp2wAmRft0mIM = 16'sb0000000000000000; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : j2gHN9roTaQcXLtCUWIL9F if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin k9BY0fd7LFxuaZBtnq2NstC[0] <= 16'sb0000000000000000; k9BY0fd7LFxuaZBtnq2NstC[1] <= 16'sb0000000000000000; k9BY0fd7LFxuaZBtnq2NstC[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin k9BY0fd7LFxuaZBtnq2NstC[0] <= 16'sb0000000000000000; k9BY0fd7LFxuaZBtnq2NstC[1] <= 16'sb0000000000000000; k9BY0fd7LFxuaZBtnq2NstC[2] <= 16'sb0000000000000000; end else begin k9BY0fd7LFxuaZBtnq2NstC[0] <= mTZgUkGw3710r8TqEV6XWF[0]; k9BY0fd7LFxuaZBtnq2NstC[1] <= mTZgUkGw3710r8TqEV6XWF[1]; k9BY0fd7LFxuaZBtnq2NstC[2] <= mTZgUkGw3710r8TqEV6XWF[2]; end end end assign sueXASR1jeFcZWA77t3pGH = k9BY0fd7LFxuaZBtnq2NstC[2]; assign mTZgUkGw3710r8TqEV6XWF[0] = KD169OZrhp2wAmRft0mIM; assign mTZgUkGw3710r8TqEV6XWF[1] = k9BY0fd7LFxuaZBtnq2NstC[0]; assign mTZgUkGw3710r8TqEV6XWF[2] = k9BY0fd7LFxuaZBtnq2NstC[1]; DoB23Fa4uAIKH4YzWRxQJC qlkqShI2B6dsvULpxRGpgG (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .RclzV3Jlkk5FKKnL0G6JcF(RclzV3Jlkk5FKKnL0G6JcF), .sueXASR1jeFcZWA77t3pGH(sueXASR1jeFcZWA77t3pGH), .JdpDaA8gpSp0rE35OGZkGE(JdpDaA8gpSp0rE35OGZkGE), .u5bboUjXYRZBbt1duYbKTG(u5bboUjXYRZBbt1duYbKTG), .mir92X5UlUGvLQSXmCuq9(mir92X5UlUGvLQSXmCuq9), .hOMBB3qOa4Z6E9dukDYA0F(hOMBB3qOa4Z6E9dukDYA0F), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .d41CUYvsIlUzO1gIRNNShD(d41CUYvsIlUzO1gIRNNShD), .QLKtWBpH0VjEHhv0F6cEGD(QLKtWBpH0VjEHhv0F6cEGD) ); ZKzJfveV1YombAboWD3IdD JvzDhpwb7aUlHKaT7fPbLF (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .d41CUYvsIlUzO1gIRNNShD(d41CUYvsIlUzO1gIRNNShD), .QLKtWBpH0VjEHhv0F6cEGD(QLKtWBpH0VjEHhv0F6cEGD), .c070CKvbOwMMYffRzNpxjuG(c070CKvbOwMMYffRzNpxjuG), .BZMbpSF4BAilhRWeHczrfC(BZMbpSF4BAilhRWeHczrfC), .Ax88y9n8GnrKjg0yG0FKzE(Ax88y9n8GnrKjg0yG0FKzE), .CosmSfOlF9hl7OPB7KnKvB(CosmSfOlF9hl7OPB7KnKvB), .rFrTP2XEQaUmbjytbnblxB(rFrTP2XEQaUmbjytbnblxB), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .LHOKWpKrWmWJXxxXqAj0TH(LHOKWpKrWmWJXxxXqAj0TH), .u9UFtyHKgbvGPJXvb5sSmF(u9UFtyHKgbvGPJXvb5sSmF) ); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : eVDXDpbSTruDFXBM6ygPaB if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin k8gGlV5iKkuIBPqjsMS5KF[0] <= 16'sb0000000000000000; k8gGlV5iKkuIBPqjsMS5KF[1] <= 16'sb0000000000000000; k8gGlV5iKkuIBPqjsMS5KF[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin k8gGlV5iKkuIBPqjsMS5KF[0] <= 16'sb0000000000000000; k8gGlV5iKkuIBPqjsMS5KF[1] <= 16'sb0000000000000000; k8gGlV5iKkuIBPqjsMS5KF[2] <= 16'sb0000000000000000; end else begin k8gGlV5iKkuIBPqjsMS5KF[0] <= jVudy6rBy3pL4AAajihjvH[0]; k8gGlV5iKkuIBPqjsMS5KF[1] <= jVudy6rBy3pL4AAajihjvH[1]; k8gGlV5iKkuIBPqjsMS5KF[2] <= jVudy6rBy3pL4AAajihjvH[2]; end end end assign DbYwoM2JCYD9mwcRRKmb6G = k8gGlV5iKkuIBPqjsMS5KF[2]; assign jVudy6rBy3pL4AAajihjvH[0] = LHOKWpKrWmWJXxxXqAj0TH; assign jVudy6rBy3pL4AAajihjvH[1] = k8gGlV5iKkuIBPqjsMS5KF[0]; assign jVudy6rBy3pL4AAajihjvH[2] = k8gGlV5iKkuIBPqjsMS5KF[1]; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : a2bprYW6bhaVvTUhwUfmVQF if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin x9EdsEkQtjpM4w517iGHzC[0] <= 16'sb0000000000000000; x9EdsEkQtjpM4w517iGHzC[1] <= 16'sb0000000000000000; x9EdsEkQtjpM4w517iGHzC[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin x9EdsEkQtjpM4w517iGHzC[0] <= 16'sb0000000000000000; x9EdsEkQtjpM4w517iGHzC[1] <= 16'sb0000000000000000; x9EdsEkQtjpM4w517iGHzC[2] <= 16'sb0000000000000000; end else begin x9EdsEkQtjpM4w517iGHzC[0] <= tnuZKwedoQlWAtzBo6aIZB[0]; x9EdsEkQtjpM4w517iGHzC[1] <= tnuZKwedoQlWAtzBo6aIZB[1]; x9EdsEkQtjpM4w517iGHzC[2] <= tnuZKwedoQlWAtzBo6aIZB[2]; end end end assign WbySmFpEqdJe6nrpd6KgG = x9EdsEkQtjpM4w517iGHzC[2]; assign tnuZKwedoQlWAtzBo6aIZB[0] = u9UFtyHKgbvGPJXvb5sSmF; assign tnuZKwedoQlWAtzBo6aIZB[1] = x9EdsEkQtjpM4w517iGHzC[0]; assign tnuZKwedoQlWAtzBo6aIZB[2] = x9EdsEkQtjpM4w517iGHzC[1]; CWClvr8Mr00imcOxbxkVdE FYP2YP6G2rKauewwkvNbYC (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .b93Ikbo3dw8VtPD6KcPt3C(b93Ikbo3dw8VtPD6KcPt3C), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .i4y6Td18s9Zr0JbepLQtjC(i4y6Td18s9Zr0JbepLQtjC), .k3FlrGNoOUOhUgHDIDYGouE(k3FlrGNoOUOhUgHDIDYGouE) ); tCsMfmFmjTaltCEQMQbsYD w92e99l9cUvs69EuygaxMC (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .DbYwoM2JCYD9mwcRRKmb6G(DbYwoM2JCYD9mwcRRKmb6G), .WbySmFpEqdJe6nrpd6KgG(WbySmFpEqdJe6nrpd6KgG), .pCWATI9lTIGbmXTtLuLAGB(pCWATI9lTIGbmXTtLuLAGB), .yTf5WZbZOLm2uKwJmXk5sG(yTf5WZbZOLm2uKwJmXk5sG), .wGlnEfCkRPxniOjCaZH6XG(wGlnEfCkRPxniOjCaZH6XG), .i4y6Td18s9Zr0JbepLQtjC(i4y6Td18s9Zr0JbepLQtjC), .k3FlrGNoOUOhUgHDIDYGouE(k3FlrGNoOUOhUgHDIDYGouE), .RDvlVEJspE7WkJvNmR8a6C(RDvlVEJspE7WkJvNmR8a6C), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .t30W3eeadZl9O9RnQCafyED(t30W3eeadZl9O9RnQCafyED), .flGpcmOyc38fKmqiV5eQvF(flGpcmOyc38fKmqiV5eQvF) ); aoE6eYC95yLxVMOngSdpZC mrK9eCSSdfMzI9Yt8myOHB (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .t30W3eeadZl9O9RnQCafyED(t30W3eeadZl9O9RnQCafyED), .flGpcmOyc38fKmqiV5eQvF(flGpcmOyc38fKmqiV5eQvF), .DZol1WsbVnSldsei0SiI9E(DZol1WsbVnSldsei0SiI9E), .zqdZMmoxIs9zmnL4kATVuC(zqdZMmoxIs9zmnL4kATVuC), .a8rK4qdEuNCWHLdYbR2f8(a8rK4qdEuNCWHLdYbR2f8), .O6TgnxqnGk692qEmnZQFTC(O6TgnxqnGk692qEmnZQFTC), .XfCDnggI1Y1qaMzSOLL0TD(XfCDnggI1Y1qaMzSOLL0TD), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .CBqrXFTnHQDD2JNQjTxpkH(CBqrXFTnHQDD2JNQjTxpkH), .dYQ3fSOENqw4ZimOQmMMTH(dYQ3fSOENqw4ZimOQmMMTH) ); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : RfFhiu7TcZArCuQWZZoVsB if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin KmuHj4FutgT59Q7oCiggpD[0] <= 16'sb0000000000000000; KmuHj4FutgT59Q7oCiggpD[1] <= 16'sb0000000000000000; KmuHj4FutgT59Q7oCiggpD[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin KmuHj4FutgT59Q7oCiggpD[0] <= 16'sb0000000000000000; KmuHj4FutgT59Q7oCiggpD[1] <= 16'sb0000000000000000; KmuHj4FutgT59Q7oCiggpD[2] <= 16'sb0000000000000000; end else begin KmuHj4FutgT59Q7oCiggpD[0] <= UFFCUGMTW5jYs8JEV3j3KC[0]; KmuHj4FutgT59Q7oCiggpD[1] <= UFFCUGMTW5jYs8JEV3j3KC[1]; KmuHj4FutgT59Q7oCiggpD[2] <= UFFCUGMTW5jYs8JEV3j3KC[2]; end end end assign lSTAIQPANZYVi9u1bQJbfC = KmuHj4FutgT59Q7oCiggpD[2]; assign UFFCUGMTW5jYs8JEV3j3KC[0] = CBqrXFTnHQDD2JNQjTxpkH; assign UFFCUGMTW5jYs8JEV3j3KC[1] = KmuHj4FutgT59Q7oCiggpD[0]; assign UFFCUGMTW5jYs8JEV3j3KC[2] = KmuHj4FutgT59Q7oCiggpD[1]; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : owLoaMKUokO7uUwJJovpJE if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin appAG8sqUT59wY8ObKEssF[0] <= 16'sb0000000000000000; appAG8sqUT59wY8ObKEssF[1] <= 16'sb0000000000000000; appAG8sqUT59wY8ObKEssF[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin appAG8sqUT59wY8ObKEssF[0] <= 16'sb0000000000000000; appAG8sqUT59wY8ObKEssF[1] <= 16'sb0000000000000000; appAG8sqUT59wY8ObKEssF[2] <= 16'sb0000000000000000; end else begin appAG8sqUT59wY8ObKEssF[0] <= d21AAbScpxqwLWzuGxj8ajB[0]; appAG8sqUT59wY8ObKEssF[1] <= d21AAbScpxqwLWzuGxj8ajB[1]; appAG8sqUT59wY8ObKEssF[2] <= d21AAbScpxqwLWzuGxj8ajB[2]; end end end assign hh7M8p6TyfjHKgE0YxcN3 = appAG8sqUT59wY8ObKEssF[2]; assign d21AAbScpxqwLWzuGxj8ajB[0] = dYQ3fSOENqw4ZimOQmMMTH; assign d21AAbScpxqwLWzuGxj8ajB[1] = appAG8sqUT59wY8ObKEssF[0]; assign d21AAbScpxqwLWzuGxj8ajB[2] = appAG8sqUT59wY8ObKEssF[1]; v1FZ9BAyYkzKAQiHSjAsZyC k9LBugZcaE827GA1WMmAUmF (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .NMWfejbHi1tIjFkylFWDkC(NMWfejbHi1tIjFkylFWDkC), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .FB6nKajjqrTT1538hBpQ9C(FB6nKajjqrTT1538hBpQ9C), .XcmpMS0nhYnUzTPGBkEmmF(XcmpMS0nhYnUzTPGBkEmmF) ); r8TsfnOtUTBk35ooa4HDQAD rwgHjaAP6nzyxxSYcq7lpF (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .lSTAIQPANZYVi9u1bQJbfC(lSTAIQPANZYVi9u1bQJbfC), .hh7M8p6TyfjHKgE0YxcN3(hh7M8p6TyfjHKgE0YxcN3), .v6PtMRDEb2KzMpzXWCSiwkB(v6PtMRDEb2KzMpzXWCSiwkB), .u6oVvmCf0f079jLPodlV5B(u6oVvmCf0f079jLPodlV5B), .qv4pS1KBm1VYTuOTZHo04F(qv4pS1KBm1VYTuOTZHo04F), .FB6nKajjqrTT1538hBpQ9C(FB6nKajjqrTT1538hBpQ9C), .XcmpMS0nhYnUzTPGBkEmmF(XcmpMS0nhYnUzTPGBkEmmF), .LSv5mOYTPLq5vaIpiVTypC(LSv5mOYTPLq5vaIpiVTypC), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .OAkG388GVoqfAFfrsC3Z3(OAkG388GVoqfAFfrsC3Z3), .DP58bSOk4VSBFH6tnqlVTH(DP58bSOk4VSBFH6tnqlVTH) ); IT7y3HrJPu7teNsd6CIHy qain7iDZFbUFjqzZeJib6E (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .OAkG388GVoqfAFfrsC3Z3(OAkG388GVoqfAFfrsC3Z3), .DP58bSOk4VSBFH6tnqlVTH(DP58bSOk4VSBFH6tnqlVTH), .Ck459KQ1C8vRbine3lrkt(Ck459KQ1C8vRbine3lrkt), .MCqIdNMOB0Mg1cefHLMjpH(MCqIdNMOB0Mg1cefHLMjpH), .j41GwwL8b9NI9l6ZScQ1PbG(j41GwwL8b9NI9l6ZScQ1PbG), .i8H7HzN3cvjFks6MZ5qaqF(i8H7HzN3cvjFks6MZ5qaqF), .SAcShGLK2YZQrWHGqGVvjD(SAcShGLK2YZQrWHGqGVvjD), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .oEtRmwXRZkMV2JHZdumYM(oEtRmwXRZkMV2JHZdumYM), .ABAJKgUy1j1LH4rwhRtEnG(ABAJKgUy1j1LH4rwhRtEnG) ); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : YKhHebQtfFPtGJB8AN9NfC if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin pISZVQJtPY1M87J4LAx1MB[0] <= 16'sb0000000000000000; pISZVQJtPY1M87J4LAx1MB[1] <= 16'sb0000000000000000; pISZVQJtPY1M87J4LAx1MB[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin pISZVQJtPY1M87J4LAx1MB[0] <= 16'sb0000000000000000; pISZVQJtPY1M87J4LAx1MB[1] <= 16'sb0000000000000000; pISZVQJtPY1M87J4LAx1MB[2] <= 16'sb0000000000000000; end else begin pISZVQJtPY1M87J4LAx1MB[0] <= EwyTeOtw0Znxv6WUZIsKtH[0]; pISZVQJtPY1M87J4LAx1MB[1] <= EwyTeOtw0Znxv6WUZIsKtH[1]; pISZVQJtPY1M87J4LAx1MB[2] <= EwyTeOtw0Znxv6WUZIsKtH[2]; end end end assign OTz07QnhICRdmhJUaCsjDD = pISZVQJtPY1M87J4LAx1MB[2]; assign EwyTeOtw0Znxv6WUZIsKtH[0] = oEtRmwXRZkMV2JHZdumYM; assign EwyTeOtw0Znxv6WUZIsKtH[1] = pISZVQJtPY1M87J4LAx1MB[0]; assign EwyTeOtw0Znxv6WUZIsKtH[2] = pISZVQJtPY1M87J4LAx1MB[1]; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : R02gF8dBxGuXtqNBiytOBD if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin ufyCKBsm7ZcDMoHa9lVT8B[0] <= 16'sb0000000000000000; ufyCKBsm7ZcDMoHa9lVT8B[1] <= 16'sb0000000000000000; ufyCKBsm7ZcDMoHa9lVT8B[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin ufyCKBsm7ZcDMoHa9lVT8B[0] <= 16'sb0000000000000000; ufyCKBsm7ZcDMoHa9lVT8B[1] <= 16'sb0000000000000000; ufyCKBsm7ZcDMoHa9lVT8B[2] <= 16'sb0000000000000000; end else begin ufyCKBsm7ZcDMoHa9lVT8B[0] <= lc0FzXjU6ruJOOuwpT5PQ[0]; ufyCKBsm7ZcDMoHa9lVT8B[1] <= lc0FzXjU6ruJOOuwpT5PQ[1]; ufyCKBsm7ZcDMoHa9lVT8B[2] <= lc0FzXjU6ruJOOuwpT5PQ[2]; end end end assign jnRu1hLACcXOUmEbgPMwFH = ufyCKBsm7ZcDMoHa9lVT8B[2]; assign lc0FzXjU6ruJOOuwpT5PQ[0] = ABAJKgUy1j1LH4rwhRtEnG; assign lc0FzXjU6ruJOOuwpT5PQ[1] = ufyCKBsm7ZcDMoHa9lVT8B[0]; assign lc0FzXjU6ruJOOuwpT5PQ[2] = ufyCKBsm7ZcDMoHa9lVT8B[1]; ZVnVljYRwutZ211zPnsNmD bQVBAnxXJylfCrtgM5vSPE (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .mm30CTneMiOZJcmmoHkb2D(mm30CTneMiOZJcmmoHkb2D), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .NQfJJVPm8CcUv19grKEsZB(NQfJJVPm8CcUv19grKEsZB), .k67mERxT6pCrtuCZzqKAJD(k67mERxT6pCrtuCZzqKAJD) ); EDdmCjHV1lGAjBmFyUBFmB i7dnMCtdoD6bNq2cmT7P1E (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .OTz07QnhICRdmhJUaCsjDD(OTz07QnhICRdmhJUaCsjDD), .jnRu1hLACcXOUmEbgPMwFH(jnRu1hLACcXOUmEbgPMwFH), .l9QVSAqS6jsMaipvGnosLD(l9QVSAqS6jsMaipvGnosLD), .g1oJwDFAtNAcPvLahTlMEB(g1oJwDFAtNAcPvLahTlMEB), .wf5f4XnltnQYt1bEDWEp0F(wf5f4XnltnQYt1bEDWEp0F), .NQfJJVPm8CcUv19grKEsZB(NQfJJVPm8CcUv19grKEsZB), .k67mERxT6pCrtuCZzqKAJD(k67mERxT6pCrtuCZzqKAJD), .Q7D2KKVRLkwEPktPhyCkSD(Q7D2KKVRLkwEPktPhyCkSD), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .lZzpoGgoYZNYjthSDnLuPH(lZzpoGgoYZNYjthSDnLuPH), .R8WEgTosuCMkRIvxet0i5D(R8WEgTosuCMkRIvxet0i5D) ); uORIqLwjUCOEz15zmk6d4C gAoRepPamcDhvSXs2STBZ (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .lZzpoGgoYZNYjthSDnLuPH(lZzpoGgoYZNYjthSDnLuPH), .R8WEgTosuCMkRIvxet0i5D(R8WEgTosuCMkRIvxet0i5D), .QWAACQosHJOUrDgm1wJeoG(QWAACQosHJOUrDgm1wJeoG), .WgU2KCxd1j6m3EUCPiuf1F(WgU2KCxd1j6m3EUCPiuf1F), .y9Hu20tqKGzmg7O1xqeuAZH(y9Hu20tqKGzmg7O1xqeuAZH), .F9FfK0xrG2zVVJqYJzgfxD(F9FfK0xrG2zVVJqYJzgfxD), .xGMN0H1JXsbMHEVz1iuteB(xGMN0H1JXsbMHEVz1iuteB), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .gEaylbF1WXdCOYwXfvD4G(gEaylbF1WXdCOYwXfvD4G), .o4iXCc2GyRgQIsHmtR0i8nE(o4iXCc2GyRgQIsHmtR0i8nE) ); i4lJrvliAJeiTHUjYckKWwC zQATYzKjyddZYs5E14edv (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .NdNevEoWljk83nSbsGDU1C(NdNevEoWljk83nSbsGDU1C), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .ymBdGOgDsRajoiY9d7TZdC(ymBdGOgDsRajoiY9d7TZdC), .q8L6STCfvGEzwAAhXRTKviE(q8L6STCfvGEzwAAhXRTKviE) ); PgyJIAY0PTIwvT911tPTDC RZ1M7pkYSnFBKBsZutNghD (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .l7IYN7joqiz566PVFOWVRgE(l7IYN7joqiz566PVFOWVRgE), .WJrLCpghLrgwyLgXr83JPE(WJrLCpghLrgwyLgXr83JPE), .gEaylbF1WXdCOYwXfvD4G(gEaylbF1WXdCOYwXfvD4G), .o4iXCc2GyRgQIsHmtR0i8nE(o4iXCc2GyRgQIsHmtR0i8nE), .NdNevEoWljk83nSbsGDU1C(NdNevEoWljk83nSbsGDU1C), .ymBdGOgDsRajoiY9d7TZdC(ymBdGOgDsRajoiY9d7TZdC), .q8L6STCfvGEzwAAhXRTKviE(q8L6STCfvGEzwAAhXRTKviE), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .EnlAo7K66kKuzHIKWLmc1F(EnlAo7K66kKuzHIKWLmc1F), .ew3EeLap6s8rXmNrsqaTWH(ew3EeLap6s8rXmNrsqaTWH), .IPh1M0O3x0ioGlon72MROG(IPh1M0O3x0ioGlon72MROG), .Mt05SNCQbo0cCPNa1yEFyF(Mt05SNCQbo0cCPNa1yEFyF), .Z7ZDy0EvwvoCh1zahAqvSF(Z7ZDy0EvwvoCh1zahAqvSF) ); assign V7D51SjWfBbpNwnqW3bM8F = J5kDQbkAAS4E39jPz9JzwD; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : Fxt9eCqtG0jUXmLi6jZUvE if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin f6n0j0rIhtlF1cK7ntOhdG[0] <= 16'sb0000000000000000; f6n0j0rIhtlF1cK7ntOhdG[1] <= 16'sb0000000000000000; f6n0j0rIhtlF1cK7ntOhdG[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin f6n0j0rIhtlF1cK7ntOhdG[0] <= 16'sb0000000000000000; f6n0j0rIhtlF1cK7ntOhdG[1] <= 16'sb0000000000000000; f6n0j0rIhtlF1cK7ntOhdG[2] <= 16'sb0000000000000000; end else begin f6n0j0rIhtlF1cK7ntOhdG[0] <= f8PGb7nqRvYgidEKAnbVYCF[0]; f6n0j0rIhtlF1cK7ntOhdG[1] <= f8PGb7nqRvYgidEKAnbVYCF[1]; f6n0j0rIhtlF1cK7ntOhdG[2] <= f8PGb7nqRvYgidEKAnbVYCF[2]; end end end assign SvMbkNSHmfXxZeVeRXimM = f6n0j0rIhtlF1cK7ntOhdG[2]; assign f8PGb7nqRvYgidEKAnbVYCF[0] = V7D51SjWfBbpNwnqW3bM8F; assign f8PGb7nqRvYgidEKAnbVYCF[1] = f6n0j0rIhtlF1cK7ntOhdG[0]; assign f8PGb7nqRvYgidEKAnbVYCF[2] = f6n0j0rIhtlF1cK7ntOhdG[1]; assign a9SSaqPU7lUCu5a3eXSIsF = 16'sb0000000000000000; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : iRHyolisTvsKLxVejMexAB if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin hDe4KgCGLUE2lc3mBRHUGE[0] <= 16'sb0000000000000000; hDe4KgCGLUE2lc3mBRHUGE[1] <= 16'sb0000000000000000; hDe4KgCGLUE2lc3mBRHUGE[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin hDe4KgCGLUE2lc3mBRHUGE[0] <= 16'sb0000000000000000; hDe4KgCGLUE2lc3mBRHUGE[1] <= 16'sb0000000000000000; hDe4KgCGLUE2lc3mBRHUGE[2] <= 16'sb0000000000000000; end else begin hDe4KgCGLUE2lc3mBRHUGE[0] <= ZvqDLDMtFPbHpUtzihpbXF[0]; hDe4KgCGLUE2lc3mBRHUGE[1] <= ZvqDLDMtFPbHpUtzihpbXF[1]; hDe4KgCGLUE2lc3mBRHUGE[2] <= ZvqDLDMtFPbHpUtzihpbXF[2]; end end end assign qGH0gnrBBGm2QIOAgMsMCH = hDe4KgCGLUE2lc3mBRHUGE[2]; assign ZvqDLDMtFPbHpUtzihpbXF[0] = a9SSaqPU7lUCu5a3eXSIsF; assign ZvqDLDMtFPbHpUtzihpbXF[1] = hDe4KgCGLUE2lc3mBRHUGE[0]; assign ZvqDLDMtFPbHpUtzihpbXF[2] = hDe4KgCGLUE2lc3mBRHUGE[1]; tnJK3GkhopKNT9tFixA22D qESeGovVleC0wdJW7G4WyF (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .SvMbkNSHmfXxZeVeRXimM(SvMbkNSHmfXxZeVeRXimM), .qGH0gnrBBGm2QIOAgMsMCH(qGH0gnrBBGm2QIOAgMsMCH), .JdpDaA8gpSp0rE35OGZkGE(JdpDaA8gpSp0rE35OGZkGE), .u5bboUjXYRZBbt1duYbKTG(u5bboUjXYRZBbt1duYbKTG), .mir92X5UlUGvLQSXmCuq9(mir92X5UlUGvLQSXmCuq9), .hOMBB3qOa4Z6E9dukDYA0F(hOMBB3qOa4Z6E9dukDYA0F), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .TyWfuK18qujvo4OtMAdhe(TyWfuK18qujvo4OtMAdhe), .PoiwHvfIvYu5tuiBaljpTF(PoiwHvfIvYu5tuiBaljpTF) ); BLlulIvcVSY8PU777oEMRC o074bALxe21FtOafjH7oMH (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .TyWfuK18qujvo4OtMAdhe(TyWfuK18qujvo4OtMAdhe), .PoiwHvfIvYu5tuiBaljpTF(PoiwHvfIvYu5tuiBaljpTF), .c070CKvbOwMMYffRzNpxjuG(c070CKvbOwMMYffRzNpxjuG), .BZMbpSF4BAilhRWeHczrfC(BZMbpSF4BAilhRWeHczrfC), .Ax88y9n8GnrKjg0yG0FKzE(Ax88y9n8GnrKjg0yG0FKzE), .CosmSfOlF9hl7OPB7KnKvB(CosmSfOlF9hl7OPB7KnKvB), .rFrTP2XEQaUmbjytbnblxB(rFrTP2XEQaUmbjytbnblxB), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .WdhKnVKybfbzc7shj6T5ID(WdhKnVKybfbzc7shj6T5ID), .Z8VgU0v1VN5pqpZolA5AtF(Z8VgU0v1VN5pqpZolA5AtF) ); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : e6AZe9KIcZJURxtpakQhtqG if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin I3TwcvTY4hEZBUKyNKGQYH[0] <= 16'sb0000000000000000; I3TwcvTY4hEZBUKyNKGQYH[1] <= 16'sb0000000000000000; I3TwcvTY4hEZBUKyNKGQYH[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin I3TwcvTY4hEZBUKyNKGQYH[0] <= 16'sb0000000000000000; I3TwcvTY4hEZBUKyNKGQYH[1] <= 16'sb0000000000000000; I3TwcvTY4hEZBUKyNKGQYH[2] <= 16'sb0000000000000000; end else begin I3TwcvTY4hEZBUKyNKGQYH[0] <= ltutKZEJ3uAsYBtveZfxN[0]; I3TwcvTY4hEZBUKyNKGQYH[1] <= ltutKZEJ3uAsYBtveZfxN[1]; I3TwcvTY4hEZBUKyNKGQYH[2] <= ltutKZEJ3uAsYBtveZfxN[2]; end end end assign risZnLFYvPBrH1cy6dfHMF = I3TwcvTY4hEZBUKyNKGQYH[2]; assign ltutKZEJ3uAsYBtveZfxN[0] = WdhKnVKybfbzc7shj6T5ID; assign ltutKZEJ3uAsYBtveZfxN[1] = I3TwcvTY4hEZBUKyNKGQYH[0]; assign ltutKZEJ3uAsYBtveZfxN[2] = I3TwcvTY4hEZBUKyNKGQYH[1]; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : y8LVueovJyghRSuIm8a5QH if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin h41dWYc0X3ZAsDk44FMtsTD[0] <= 16'sb0000000000000000; h41dWYc0X3ZAsDk44FMtsTD[1] <= 16'sb0000000000000000; h41dWYc0X3ZAsDk44FMtsTD[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin h41dWYc0X3ZAsDk44FMtsTD[0] <= 16'sb0000000000000000; h41dWYc0X3ZAsDk44FMtsTD[1] <= 16'sb0000000000000000; h41dWYc0X3ZAsDk44FMtsTD[2] <= 16'sb0000000000000000; end else begin h41dWYc0X3ZAsDk44FMtsTD[0] <= kZIaatjtNR5S1owTPfmSI[0]; h41dWYc0X3ZAsDk44FMtsTD[1] <= kZIaatjtNR5S1owTPfmSI[1]; h41dWYc0X3ZAsDk44FMtsTD[2] <= kZIaatjtNR5S1owTPfmSI[2]; end end end assign y3mUIhc5hpdbI6gB0Klf3MH = h41dWYc0X3ZAsDk44FMtsTD[2]; assign kZIaatjtNR5S1owTPfmSI[0] = Z8VgU0v1VN5pqpZolA5AtF; assign kZIaatjtNR5S1owTPfmSI[1] = h41dWYc0X3ZAsDk44FMtsTD[0]; assign kZIaatjtNR5S1owTPfmSI[2] = h41dWYc0X3ZAsDk44FMtsTD[1]; cN8kZ5KZqHVjQmLZPPEnXH rbo4XnEDAmRflkh99n2moB (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .b93Ikbo3dw8VtPD6KcPt3C(b93Ikbo3dw8VtPD6KcPt3C), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .UlGc2PVtJa9BNobxUHDxSG(UlGc2PVtJa9BNobxUHDxSG), .pdTCH0gTlgy9qR74rtvuBE(pdTCH0gTlgy9qR74rtvuBE) ); f25aX5QlpO938C34Yy3CBdC ryVcsu5GzuSm41uBLdn2YE (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .risZnLFYvPBrH1cy6dfHMF(risZnLFYvPBrH1cy6dfHMF), .y3mUIhc5hpdbI6gB0Klf3MH(y3mUIhc5hpdbI6gB0Klf3MH), .pCWATI9lTIGbmXTtLuLAGB(pCWATI9lTIGbmXTtLuLAGB), .yTf5WZbZOLm2uKwJmXk5sG(yTf5WZbZOLm2uKwJmXk5sG), .wGlnEfCkRPxniOjCaZH6XG(wGlnEfCkRPxniOjCaZH6XG), .UlGc2PVtJa9BNobxUHDxSG(UlGc2PVtJa9BNobxUHDxSG), .pdTCH0gTlgy9qR74rtvuBE(pdTCH0gTlgy9qR74rtvuBE), .RDvlVEJspE7WkJvNmR8a6C(RDvlVEJspE7WkJvNmR8a6C), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .msLJn85q5aDnigXPSLnA9F(msLJn85q5aDnigXPSLnA9F), .s8tbEDkTdSLkOXc5hVDArH(s8tbEDkTdSLkOXc5hVDArH) ); LeezLu8utZvbs8zm8S97TD ef4GM1uMXwhosxoRlEdZMF (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .msLJn85q5aDnigXPSLnA9F(msLJn85q5aDnigXPSLnA9F), .s8tbEDkTdSLkOXc5hVDArH(s8tbEDkTdSLkOXc5hVDArH), .DZol1WsbVnSldsei0SiI9E(DZol1WsbVnSldsei0SiI9E), .zqdZMmoxIs9zmnL4kATVuC(zqdZMmoxIs9zmnL4kATVuC), .a8rK4qdEuNCWHLdYbR2f8(a8rK4qdEuNCWHLdYbR2f8), .O6TgnxqnGk692qEmnZQFTC(O6TgnxqnGk692qEmnZQFTC), .XfCDnggI1Y1qaMzSOLL0TD(XfCDnggI1Y1qaMzSOLL0TD), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .ACHpp43jQbQJO4HdGlLQ0B(ACHpp43jQbQJO4HdGlLQ0B), .BJNXQzaMpa7r8LYTHlOrBD(BJNXQzaMpa7r8LYTHlOrBD) ); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : Yera4SjAVuKG7TjeL0xum if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin UbhppxZFtuRiGSMYxgMT2F[0] <= 16'sb0000000000000000; UbhppxZFtuRiGSMYxgMT2F[1] <= 16'sb0000000000000000; UbhppxZFtuRiGSMYxgMT2F[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin UbhppxZFtuRiGSMYxgMT2F[0] <= 16'sb0000000000000000; UbhppxZFtuRiGSMYxgMT2F[1] <= 16'sb0000000000000000; UbhppxZFtuRiGSMYxgMT2F[2] <= 16'sb0000000000000000; end else begin UbhppxZFtuRiGSMYxgMT2F[0] <= rk6XtqxIQmYnoKIvpO9PNH[0]; UbhppxZFtuRiGSMYxgMT2F[1] <= rk6XtqxIQmYnoKIvpO9PNH[1]; UbhppxZFtuRiGSMYxgMT2F[2] <= rk6XtqxIQmYnoKIvpO9PNH[2]; end end end assign BXAaMHpKzPpYZGFRqoevNE = UbhppxZFtuRiGSMYxgMT2F[2]; assign rk6XtqxIQmYnoKIvpO9PNH[0] = ACHpp43jQbQJO4HdGlLQ0B; assign rk6XtqxIQmYnoKIvpO9PNH[1] = UbhppxZFtuRiGSMYxgMT2F[0]; assign rk6XtqxIQmYnoKIvpO9PNH[2] = UbhppxZFtuRiGSMYxgMT2F[1]; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : MplkH2AOPP4uw14V7wrk3B if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin TGSVeodh4aSh5YMUFsJBpF[0] <= 16'sb0000000000000000; TGSVeodh4aSh5YMUFsJBpF[1] <= 16'sb0000000000000000; TGSVeodh4aSh5YMUFsJBpF[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin TGSVeodh4aSh5YMUFsJBpF[0] <= 16'sb0000000000000000; TGSVeodh4aSh5YMUFsJBpF[1] <= 16'sb0000000000000000; TGSVeodh4aSh5YMUFsJBpF[2] <= 16'sb0000000000000000; end else begin TGSVeodh4aSh5YMUFsJBpF[0] <= pKwMCjbBuwX4wlYrJtZeqH[0]; TGSVeodh4aSh5YMUFsJBpF[1] <= pKwMCjbBuwX4wlYrJtZeqH[1]; TGSVeodh4aSh5YMUFsJBpF[2] <= pKwMCjbBuwX4wlYrJtZeqH[2]; end end end assign czP63K90EaJdtsY9EHZ30D = TGSVeodh4aSh5YMUFsJBpF[2]; assign pKwMCjbBuwX4wlYrJtZeqH[0] = BJNXQzaMpa7r8LYTHlOrBD; assign pKwMCjbBuwX4wlYrJtZeqH[1] = TGSVeodh4aSh5YMUFsJBpF[0]; assign pKwMCjbBuwX4wlYrJtZeqH[2] = TGSVeodh4aSh5YMUFsJBpF[1]; ZQUjbjy2Q8cHV0ObA5D1WC rq8qvMxzcI3hsMYdni7iCG (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .NMWfejbHi1tIjFkylFWDkC(NMWfejbHi1tIjFkylFWDkC), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .mxtJaiWQH83FcZ66WqnMiH(mxtJaiWQH83FcZ66WqnMiH), .MtlWbaE0z2xTCIy368PlWF(MtlWbaE0z2xTCIy368PlWF) ); esVSS9XtBKzKANShQjPOMH NueGwXUbsNsksA8LXNYmz (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .BXAaMHpKzPpYZGFRqoevNE(BXAaMHpKzPpYZGFRqoevNE), .czP63K90EaJdtsY9EHZ30D(czP63K90EaJdtsY9EHZ30D), .v6PtMRDEb2KzMpzXWCSiwkB(v6PtMRDEb2KzMpzXWCSiwkB), .u6oVvmCf0f079jLPodlV5B(u6oVvmCf0f079jLPodlV5B), .qv4pS1KBm1VYTuOTZHo04F(qv4pS1KBm1VYTuOTZHo04F), .mxtJaiWQH83FcZ66WqnMiH(mxtJaiWQH83FcZ66WqnMiH), .MtlWbaE0z2xTCIy368PlWF(MtlWbaE0z2xTCIy368PlWF), .LSv5mOYTPLq5vaIpiVTypC(LSv5mOYTPLq5vaIpiVTypC), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .Sek0doTmbyRuabtHW5JKgH(Sek0doTmbyRuabtHW5JKgH), .h4q2yYljVPy2UhMxEpHXfqG(h4q2yYljVPy2UhMxEpHXfqG) ); iIsgOdVtTXcPw31pLI8fkC yJxVRtqjhNAc0K7yzwOlqF (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .Sek0doTmbyRuabtHW5JKgH(Sek0doTmbyRuabtHW5JKgH), .h4q2yYljVPy2UhMxEpHXfqG(h4q2yYljVPy2UhMxEpHXfqG), .Ck459KQ1C8vRbine3lrkt(Ck459KQ1C8vRbine3lrkt), .MCqIdNMOB0Mg1cefHLMjpH(MCqIdNMOB0Mg1cefHLMjpH), .j41GwwL8b9NI9l6ZScQ1PbG(j41GwwL8b9NI9l6ZScQ1PbG), .i8H7HzN3cvjFks6MZ5qaqF(i8H7HzN3cvjFks6MZ5qaqF), .SAcShGLK2YZQrWHGqGVvjD(SAcShGLK2YZQrWHGqGVvjD), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .Ni5CWVNOepdNWeLhPbktyC(Ni5CWVNOepdNWeLhPbktyC), .oC9IZ8suhbNZiMMpUwYFZE(oC9IZ8suhbNZiMMpUwYFZE) ); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : QkTsAMX2ysQgjvkiAUs2oC if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin t1XxIWfdmuGYgMJ14AA5aoF[0] <= 16'sb0000000000000000; t1XxIWfdmuGYgMJ14AA5aoF[1] <= 16'sb0000000000000000; t1XxIWfdmuGYgMJ14AA5aoF[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin t1XxIWfdmuGYgMJ14AA5aoF[0] <= 16'sb0000000000000000; t1XxIWfdmuGYgMJ14AA5aoF[1] <= 16'sb0000000000000000; t1XxIWfdmuGYgMJ14AA5aoF[2] <= 16'sb0000000000000000; end else begin t1XxIWfdmuGYgMJ14AA5aoF[0] <= Ed8ZUSDNSkOaxlQSyerJMG[0]; t1XxIWfdmuGYgMJ14AA5aoF[1] <= Ed8ZUSDNSkOaxlQSyerJMG[1]; t1XxIWfdmuGYgMJ14AA5aoF[2] <= Ed8ZUSDNSkOaxlQSyerJMG[2]; end end end assign lTYYhj3P59f6KeSXhObJAE = t1XxIWfdmuGYgMJ14AA5aoF[2]; assign Ed8ZUSDNSkOaxlQSyerJMG[0] = Ni5CWVNOepdNWeLhPbktyC; assign Ed8ZUSDNSkOaxlQSyerJMG[1] = t1XxIWfdmuGYgMJ14AA5aoF[0]; assign Ed8ZUSDNSkOaxlQSyerJMG[2] = t1XxIWfdmuGYgMJ14AA5aoF[1]; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : EUqbtBsMjpkspgfBj9UDCG if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin u4aeKdZeegD94j2S6reFTD[0] <= 16'sb0000000000000000; u4aeKdZeegD94j2S6reFTD[1] <= 16'sb0000000000000000; u4aeKdZeegD94j2S6reFTD[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin u4aeKdZeegD94j2S6reFTD[0] <= 16'sb0000000000000000; u4aeKdZeegD94j2S6reFTD[1] <= 16'sb0000000000000000; u4aeKdZeegD94j2S6reFTD[2] <= 16'sb0000000000000000; end else begin u4aeKdZeegD94j2S6reFTD[0] <= UAnK8iuwkF7gLvWzaOGeMF[0]; u4aeKdZeegD94j2S6reFTD[1] <= UAnK8iuwkF7gLvWzaOGeMF[1]; u4aeKdZeegD94j2S6reFTD[2] <= UAnK8iuwkF7gLvWzaOGeMF[2]; end end end assign WawYOEnpsrkHlANz6YaiLG = u4aeKdZeegD94j2S6reFTD[2]; assign UAnK8iuwkF7gLvWzaOGeMF[0] = oC9IZ8suhbNZiMMpUwYFZE; assign UAnK8iuwkF7gLvWzaOGeMF[1] = u4aeKdZeegD94j2S6reFTD[0]; assign UAnK8iuwkF7gLvWzaOGeMF[2] = u4aeKdZeegD94j2S6reFTD[1]; BtkjFhnzg4iAVqQUj55ZBC F90JVXWaKZWqArerfGE6dF (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .mm30CTneMiOZJcmmoHkb2D(mm30CTneMiOZJcmmoHkb2D), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .UwIsRF8C7ejj45D9sxKqgB(UwIsRF8C7ejj45D9sxKqgB), .XVoYQfnVFtlWlmN3BG5OI(XVoYQfnVFtlWlmN3BG5OI) ); wp1dPKRLgUiS6J0V5WND0F WlJfdhgnvLpsOOjWRR7g9G (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .lTYYhj3P59f6KeSXhObJAE(lTYYhj3P59f6KeSXhObJAE), .WawYOEnpsrkHlANz6YaiLG(WawYOEnpsrkHlANz6YaiLG), .l9QVSAqS6jsMaipvGnosLD(l9QVSAqS6jsMaipvGnosLD), .g1oJwDFAtNAcPvLahTlMEB(g1oJwDFAtNAcPvLahTlMEB), .wf5f4XnltnQYt1bEDWEp0F(wf5f4XnltnQYt1bEDWEp0F), .UwIsRF8C7ejj45D9sxKqgB(UwIsRF8C7ejj45D9sxKqgB), .XVoYQfnVFtlWlmN3BG5OI(XVoYQfnVFtlWlmN3BG5OI), .Q7D2KKVRLkwEPktPhyCkSD(Q7D2KKVRLkwEPktPhyCkSD), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .BSsYK6f7nJDXvl3FdklrNE(BSsYK6f7nJDXvl3FdklrNE), .gGYwPRSrxVg8T85ahN6sK(gGYwPRSrxVg8T85ahN6sK) ); lfocSe94ipPcZI7FbavOlD l4bLRF5grfDEM8f7fPxdIB (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .BSsYK6f7nJDXvl3FdklrNE(BSsYK6f7nJDXvl3FdklrNE), .gGYwPRSrxVg8T85ahN6sK(gGYwPRSrxVg8T85ahN6sK), .QWAACQosHJOUrDgm1wJeoG(QWAACQosHJOUrDgm1wJeoG), .WgU2KCxd1j6m3EUCPiuf1F(WgU2KCxd1j6m3EUCPiuf1F), .y9Hu20tqKGzmg7O1xqeuAZH(y9Hu20tqKGzmg7O1xqeuAZH), .F9FfK0xrG2zVVJqYJzgfxD(F9FfK0xrG2zVVJqYJzgfxD), .xGMN0H1JXsbMHEVz1iuteB(xGMN0H1JXsbMHEVz1iuteB), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .S6Ue4SxCiz8dBHTO2guOUE(S6Ue4SxCiz8dBHTO2guOUE), .POhLmCr6emegQDte8TzyQ(POhLmCr6emegQDte8TzyQ) ); assign CyGvS8xQz9obtGAMlB4YwE = PVNB5uj77jMa2DXz4vJtIH; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : Hh9lAYLJ6NfTidi3vB0TOE if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin G3KM4o4fYtZmkhM463zMWE[0] <= 16'sb0000000000000000; G3KM4o4fYtZmkhM463zMWE[1] <= 16'sb0000000000000000; G3KM4o4fYtZmkhM463zMWE[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin G3KM4o4fYtZmkhM463zMWE[0] <= 16'sb0000000000000000; G3KM4o4fYtZmkhM463zMWE[1] <= 16'sb0000000000000000; G3KM4o4fYtZmkhM463zMWE[2] <= 16'sb0000000000000000; end else begin G3KM4o4fYtZmkhM463zMWE[0] <= drYAp2dAOmGqd7jeMIwcRE[0]; G3KM4o4fYtZmkhM463zMWE[1] <= drYAp2dAOmGqd7jeMIwcRE[1]; G3KM4o4fYtZmkhM463zMWE[2] <= drYAp2dAOmGqd7jeMIwcRE[2]; end end end assign TAkRd7owTLUvbZtOoRFPtC = G3KM4o4fYtZmkhM463zMWE[2]; assign drYAp2dAOmGqd7jeMIwcRE[0] = CyGvS8xQz9obtGAMlB4YwE; assign drYAp2dAOmGqd7jeMIwcRE[1] = G3KM4o4fYtZmkhM463zMWE[0]; assign drYAp2dAOmGqd7jeMIwcRE[2] = G3KM4o4fYtZmkhM463zMWE[1]; assign imE2eHPyQozGdwpwWRjBLH = 16'sb0000000000000000; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : s9hNORC8NXrLnNYPxmepXkD if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin RtR9LcVWPsx9vZqDGyBkAB[0] <= 16'sb0000000000000000; RtR9LcVWPsx9vZqDGyBkAB[1] <= 16'sb0000000000000000; RtR9LcVWPsx9vZqDGyBkAB[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin RtR9LcVWPsx9vZqDGyBkAB[0] <= 16'sb0000000000000000; RtR9LcVWPsx9vZqDGyBkAB[1] <= 16'sb0000000000000000; RtR9LcVWPsx9vZqDGyBkAB[2] <= 16'sb0000000000000000; end else begin RtR9LcVWPsx9vZqDGyBkAB[0] <= LWmwrv39ujCMpMMcrbgkHC[0]; RtR9LcVWPsx9vZqDGyBkAB[1] <= LWmwrv39ujCMpMMcrbgkHC[1]; RtR9LcVWPsx9vZqDGyBkAB[2] <= LWmwrv39ujCMpMMcrbgkHC[2]; end end end assign kj4wsLBVI5X3Usybs4WmJH = RtR9LcVWPsx9vZqDGyBkAB[2]; assign LWmwrv39ujCMpMMcrbgkHC[0] = imE2eHPyQozGdwpwWRjBLH; assign LWmwrv39ujCMpMMcrbgkHC[1] = RtR9LcVWPsx9vZqDGyBkAB[0]; assign LWmwrv39ujCMpMMcrbgkHC[2] = RtR9LcVWPsx9vZqDGyBkAB[1]; j7Pwar7D0qjQBkczNW6ZbC w34Feti8l6BGzgj9o7qjfYD (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .TAkRd7owTLUvbZtOoRFPtC(TAkRd7owTLUvbZtOoRFPtC), .kj4wsLBVI5X3Usybs4WmJH(kj4wsLBVI5X3Usybs4WmJH), .JdpDaA8gpSp0rE35OGZkGE(JdpDaA8gpSp0rE35OGZkGE), .u5bboUjXYRZBbt1duYbKTG(u5bboUjXYRZBbt1duYbKTG), .mir92X5UlUGvLQSXmCuq9(mir92X5UlUGvLQSXmCuq9), .hOMBB3qOa4Z6E9dukDYA0F(hOMBB3qOa4Z6E9dukDYA0F), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .f3NrgRvCkMfwf1E3PnKtczF(f3NrgRvCkMfwf1E3PnKtczF), .f2XZKbXdctKWPTTQYeLkBWE(f2XZKbXdctKWPTTQYeLkBWE) ); uoZ5xy8RheLCzMX3G2wpzB rRRq2JnEL8l0KURu6pY8rC (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .f3NrgRvCkMfwf1E3PnKtczF(f3NrgRvCkMfwf1E3PnKtczF), .f2XZKbXdctKWPTTQYeLkBWE(f2XZKbXdctKWPTTQYeLkBWE), .c070CKvbOwMMYffRzNpxjuG(c070CKvbOwMMYffRzNpxjuG), .BZMbpSF4BAilhRWeHczrfC(BZMbpSF4BAilhRWeHczrfC), .Ax88y9n8GnrKjg0yG0FKzE(Ax88y9n8GnrKjg0yG0FKzE), .CosmSfOlF9hl7OPB7KnKvB(CosmSfOlF9hl7OPB7KnKvB), .rFrTP2XEQaUmbjytbnblxB(rFrTP2XEQaUmbjytbnblxB), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .f6fgzNt42ufBw7e8PMAUaCB(f6fgzNt42ufBw7e8PMAUaCB), .eYtcM9qmF8eYE3uuCl3HAH(eYtcM9qmF8eYE3uuCl3HAH) ); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : g9riYEZnl9AMS1uYoZWRfJB if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin ItzBwvoI4TcHK9g7KBaUVF[0] <= 16'sb0000000000000000; ItzBwvoI4TcHK9g7KBaUVF[1] <= 16'sb0000000000000000; ItzBwvoI4TcHK9g7KBaUVF[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin ItzBwvoI4TcHK9g7KBaUVF[0] <= 16'sb0000000000000000; ItzBwvoI4TcHK9g7KBaUVF[1] <= 16'sb0000000000000000; ItzBwvoI4TcHK9g7KBaUVF[2] <= 16'sb0000000000000000; end else begin ItzBwvoI4TcHK9g7KBaUVF[0] <= fk0F6dFxBPneyImhFH4wGG[0]; ItzBwvoI4TcHK9g7KBaUVF[1] <= fk0F6dFxBPneyImhFH4wGG[1]; ItzBwvoI4TcHK9g7KBaUVF[2] <= fk0F6dFxBPneyImhFH4wGG[2]; end end end assign EiKTmNA9gqnqt6QU2ytsGF = ItzBwvoI4TcHK9g7KBaUVF[2]; assign fk0F6dFxBPneyImhFH4wGG[0] = f6fgzNt42ufBw7e8PMAUaCB; assign fk0F6dFxBPneyImhFH4wGG[1] = ItzBwvoI4TcHK9g7KBaUVF[0]; assign fk0F6dFxBPneyImhFH4wGG[2] = ItzBwvoI4TcHK9g7KBaUVF[1]; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : t21NTkKBafHvY7uJcRhS0 if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin VGCjFskQzxD0kIw7klsyNH[0] <= 16'sb0000000000000000; VGCjFskQzxD0kIw7klsyNH[1] <= 16'sb0000000000000000; VGCjFskQzxD0kIw7klsyNH[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin VGCjFskQzxD0kIw7klsyNH[0] <= 16'sb0000000000000000; VGCjFskQzxD0kIw7klsyNH[1] <= 16'sb0000000000000000; VGCjFskQzxD0kIw7klsyNH[2] <= 16'sb0000000000000000; end else begin VGCjFskQzxD0kIw7klsyNH[0] <= bsgCRrS7Pvyw5lDPgR03YH[0]; VGCjFskQzxD0kIw7klsyNH[1] <= bsgCRrS7Pvyw5lDPgR03YH[1]; VGCjFskQzxD0kIw7klsyNH[2] <= bsgCRrS7Pvyw5lDPgR03YH[2]; end end end assign i0padod73DFvzROjA4fS2o = VGCjFskQzxD0kIw7klsyNH[2]; assign bsgCRrS7Pvyw5lDPgR03YH[0] = eYtcM9qmF8eYE3uuCl3HAH; assign bsgCRrS7Pvyw5lDPgR03YH[1] = VGCjFskQzxD0kIw7klsyNH[0]; assign bsgCRrS7Pvyw5lDPgR03YH[2] = VGCjFskQzxD0kIw7klsyNH[1]; RLLhJVfo68sHjdFbtv5fcE I2TBaFHPkLkB0woW45YSD (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .b93Ikbo3dw8VtPD6KcPt3C(b93Ikbo3dw8VtPD6KcPt3C), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .mvb8xVo6CcFPFyQu3ctDE(mvb8xVo6CcFPFyQu3ctDE), .gC05dypmmuscVux3EfDHCD(gC05dypmmuscVux3EfDHCD) ); SXa0KYBbkSNWDHu83VAvL t9g2Y8fM4yk65azUUSe1E3F (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .EiKTmNA9gqnqt6QU2ytsGF(EiKTmNA9gqnqt6QU2ytsGF), .i0padod73DFvzROjA4fS2o(i0padod73DFvzROjA4fS2o), .pCWATI9lTIGbmXTtLuLAGB(pCWATI9lTIGbmXTtLuLAGB), .yTf5WZbZOLm2uKwJmXk5sG(yTf5WZbZOLm2uKwJmXk5sG), .wGlnEfCkRPxniOjCaZH6XG(wGlnEfCkRPxniOjCaZH6XG), .mvb8xVo6CcFPFyQu3ctDE(mvb8xVo6CcFPFyQu3ctDE), .gC05dypmmuscVux3EfDHCD(gC05dypmmuscVux3EfDHCD), .RDvlVEJspE7WkJvNmR8a6C(RDvlVEJspE7WkJvNmR8a6C), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .DxKKPTJNNNGcVbnDyBefdC(DxKKPTJNNNGcVbnDyBefdC), .z5IVnN9scVD1jMboeUZaZG(z5IVnN9scVD1jMboeUZaZG) ); NAZ2PhogOv6EqCFI0nhCwD bY2yqF5WO84iCOvXu7u5gH (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .DxKKPTJNNNGcVbnDyBefdC(DxKKPTJNNNGcVbnDyBefdC), .z5IVnN9scVD1jMboeUZaZG(z5IVnN9scVD1jMboeUZaZG), .DZol1WsbVnSldsei0SiI9E(DZol1WsbVnSldsei0SiI9E), .zqdZMmoxIs9zmnL4kATVuC(zqdZMmoxIs9zmnL4kATVuC), .a8rK4qdEuNCWHLdYbR2f8(a8rK4qdEuNCWHLdYbR2f8), .O6TgnxqnGk692qEmnZQFTC(O6TgnxqnGk692qEmnZQFTC), .XfCDnggI1Y1qaMzSOLL0TD(XfCDnggI1Y1qaMzSOLL0TD), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .y2F62Qir2uvIcDNjqoCgbPG(y2F62Qir2uvIcDNjqoCgbPG), .eJSHu1mAvW9BzbMy0ufWWD(eJSHu1mAvW9BzbMy0ufWWD) ); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : ocqQiwXog1G66vDmcd8fBF if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin uNvrQvd1Y0KX4XHifVskkH[0] <= 16'sb0000000000000000; uNvrQvd1Y0KX4XHifVskkH[1] <= 16'sb0000000000000000; uNvrQvd1Y0KX4XHifVskkH[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin uNvrQvd1Y0KX4XHifVskkH[0] <= 16'sb0000000000000000; uNvrQvd1Y0KX4XHifVskkH[1] <= 16'sb0000000000000000; uNvrQvd1Y0KX4XHifVskkH[2] <= 16'sb0000000000000000; end else begin uNvrQvd1Y0KX4XHifVskkH[0] <= NnZ5dINtMrF9dlFO6TR5yF[0]; uNvrQvd1Y0KX4XHifVskkH[1] <= NnZ5dINtMrF9dlFO6TR5yF[1]; uNvrQvd1Y0KX4XHifVskkH[2] <= NnZ5dINtMrF9dlFO6TR5yF[2]; end end end assign SNl44VPeKmo2uIh5zCljYE = uNvrQvd1Y0KX4XHifVskkH[2]; assign NnZ5dINtMrF9dlFO6TR5yF[0] = y2F62Qir2uvIcDNjqoCgbPG; assign NnZ5dINtMrF9dlFO6TR5yF[1] = uNvrQvd1Y0KX4XHifVskkH[0]; assign NnZ5dINtMrF9dlFO6TR5yF[2] = uNvrQvd1Y0KX4XHifVskkH[1]; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : h3NBppnMChwS5AwUtot5dF if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin keFLw9kjnIbUmEw9P3ZHlH[0] <= 16'sb0000000000000000; keFLw9kjnIbUmEw9P3ZHlH[1] <= 16'sb0000000000000000; keFLw9kjnIbUmEw9P3ZHlH[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin keFLw9kjnIbUmEw9P3ZHlH[0] <= 16'sb0000000000000000; keFLw9kjnIbUmEw9P3ZHlH[1] <= 16'sb0000000000000000; keFLw9kjnIbUmEw9P3ZHlH[2] <= 16'sb0000000000000000; end else begin keFLw9kjnIbUmEw9P3ZHlH[0] <= TdliLJ6QPHrz19i4ud5ApB[0]; keFLw9kjnIbUmEw9P3ZHlH[1] <= TdliLJ6QPHrz19i4ud5ApB[1]; keFLw9kjnIbUmEw9P3ZHlH[2] <= TdliLJ6QPHrz19i4ud5ApB[2]; end end end assign AXkTVaeFKW3Cvod76gwXK = keFLw9kjnIbUmEw9P3ZHlH[2]; assign TdliLJ6QPHrz19i4ud5ApB[0] = eJSHu1mAvW9BzbMy0ufWWD; assign TdliLJ6QPHrz19i4ud5ApB[1] = keFLw9kjnIbUmEw9P3ZHlH[0]; assign TdliLJ6QPHrz19i4ud5ApB[2] = keFLw9kjnIbUmEw9P3ZHlH[1]; MyQfGgLrTsvFkmhY4ZRirE jZAgC07ng8reotvX6puRbG (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .NMWfejbHi1tIjFkylFWDkC(NMWfejbHi1tIjFkylFWDkC), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .PV2GPYF9MTfm6A3VIE3yL(PV2GPYF9MTfm6A3VIE3yL), .VMMfdu9AIUdQe4XcwZLbSC(VMMfdu9AIUdQe4XcwZLbSC) ); JxjozggV9KBoUPlCu4g0SF x9yUjJ4dQaL4JCZ6bTAoBB (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .SNl44VPeKmo2uIh5zCljYE(SNl44VPeKmo2uIh5zCljYE), .AXkTVaeFKW3Cvod76gwXK(AXkTVaeFKW3Cvod76gwXK), .v6PtMRDEb2KzMpzXWCSiwkB(v6PtMRDEb2KzMpzXWCSiwkB), .u6oVvmCf0f079jLPodlV5B(u6oVvmCf0f079jLPodlV5B), .qv4pS1KBm1VYTuOTZHo04F(qv4pS1KBm1VYTuOTZHo04F), .PV2GPYF9MTfm6A3VIE3yL(PV2GPYF9MTfm6A3VIE3yL), .VMMfdu9AIUdQe4XcwZLbSC(VMMfdu9AIUdQe4XcwZLbSC), .LSv5mOYTPLq5vaIpiVTypC(LSv5mOYTPLq5vaIpiVTypC), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .BSA6wYLjrd40iGAxWAWPUG(BSA6wYLjrd40iGAxWAWPUG), .mVsThSJWeEPGLaZQZJ476C(mVsThSJWeEPGLaZQZJ476C) ); XumC9BzxulOwrSnrBlDCDH frmFPr2Hgpf7JABWVreFmH (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .BSA6wYLjrd40iGAxWAWPUG(BSA6wYLjrd40iGAxWAWPUG), .mVsThSJWeEPGLaZQZJ476C(mVsThSJWeEPGLaZQZJ476C), .Ck459KQ1C8vRbine3lrkt(Ck459KQ1C8vRbine3lrkt), .MCqIdNMOB0Mg1cefHLMjpH(MCqIdNMOB0Mg1cefHLMjpH), .j41GwwL8b9NI9l6ZScQ1PbG(j41GwwL8b9NI9l6ZScQ1PbG), .i8H7HzN3cvjFks6MZ5qaqF(i8H7HzN3cvjFks6MZ5qaqF), .SAcShGLK2YZQrWHGqGVvjD(SAcShGLK2YZQrWHGqGVvjD), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .Qjop49qrCNJ2RVI1tmxWK(Qjop49qrCNJ2RVI1tmxWK), .qtlf3VUxsnDXMsfKMVqqRD(qtlf3VUxsnDXMsfKMVqqRD) ); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : uFF9lWTNjcbGBQ2KohbDDF if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin a6YcmlBpfsspWdA41bdAcl[0] <= 16'sb0000000000000000; a6YcmlBpfsspWdA41bdAcl[1] <= 16'sb0000000000000000; a6YcmlBpfsspWdA41bdAcl[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin a6YcmlBpfsspWdA41bdAcl[0] <= 16'sb0000000000000000; a6YcmlBpfsspWdA41bdAcl[1] <= 16'sb0000000000000000; a6YcmlBpfsspWdA41bdAcl[2] <= 16'sb0000000000000000; end else begin a6YcmlBpfsspWdA41bdAcl[0] <= LYFiNcEj0dggwMwtkvSMMG[0]; a6YcmlBpfsspWdA41bdAcl[1] <= LYFiNcEj0dggwMwtkvSMMG[1]; a6YcmlBpfsspWdA41bdAcl[2] <= LYFiNcEj0dggwMwtkvSMMG[2]; end end end assign g86YyREiAmzs3zk0UOLK0TH = a6YcmlBpfsspWdA41bdAcl[2]; assign LYFiNcEj0dggwMwtkvSMMG[0] = Qjop49qrCNJ2RVI1tmxWK; assign LYFiNcEj0dggwMwtkvSMMG[1] = a6YcmlBpfsspWdA41bdAcl[0]; assign LYFiNcEj0dggwMwtkvSMMG[2] = a6YcmlBpfsspWdA41bdAcl[1]; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : Ptm5crw1DWlkCSU8UhL5VH if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin VLlSkvLBi8zwJgPezU50UD[0] <= 16'sb0000000000000000; VLlSkvLBi8zwJgPezU50UD[1] <= 16'sb0000000000000000; VLlSkvLBi8zwJgPezU50UD[2] <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin VLlSkvLBi8zwJgPezU50UD[0] <= 16'sb0000000000000000; VLlSkvLBi8zwJgPezU50UD[1] <= 16'sb0000000000000000; VLlSkvLBi8zwJgPezU50UD[2] <= 16'sb0000000000000000; end else begin VLlSkvLBi8zwJgPezU50UD[0] <= VLfdJwrUNkj5uYuSH99PLD[0]; VLlSkvLBi8zwJgPezU50UD[1] <= VLfdJwrUNkj5uYuSH99PLD[1]; VLlSkvLBi8zwJgPezU50UD[2] <= VLfdJwrUNkj5uYuSH99PLD[2]; end end end assign KhHmaGBWkoUJ6ybiJ9FvHH = VLlSkvLBi8zwJgPezU50UD[2]; assign VLfdJwrUNkj5uYuSH99PLD[0] = qtlf3VUxsnDXMsfKMVqqRD; assign VLfdJwrUNkj5uYuSH99PLD[1] = VLlSkvLBi8zwJgPezU50UD[0]; assign VLfdJwrUNkj5uYuSH99PLD[2] = VLlSkvLBi8zwJgPezU50UD[1]; KGrLS7nXwgj0sQ9Tard8HC iBiG4RndWj7IqE2x5Yp3eE (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .mm30CTneMiOZJcmmoHkb2D(mm30CTneMiOZJcmmoHkb2D), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .h8QlyPXT2MWg8MvvXSR0uAB(h8QlyPXT2MWg8MvvXSR0uAB), .tSs6JTBnsDJvMaRawQm6WF(tSs6JTBnsDJvMaRawQm6WF) ); Cra118G4s7bIyGNZ4oLGzB nkNufqlejWjSKGcflpnDcF (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .g86YyREiAmzs3zk0UOLK0TH(g86YyREiAmzs3zk0UOLK0TH), .KhHmaGBWkoUJ6ybiJ9FvHH(KhHmaGBWkoUJ6ybiJ9FvHH), .l9QVSAqS6jsMaipvGnosLD(l9QVSAqS6jsMaipvGnosLD), .g1oJwDFAtNAcPvLahTlMEB(g1oJwDFAtNAcPvLahTlMEB), .wf5f4XnltnQYt1bEDWEp0F(wf5f4XnltnQYt1bEDWEp0F), .h8QlyPXT2MWg8MvvXSR0uAB(h8QlyPXT2MWg8MvvXSR0uAB), .tSs6JTBnsDJvMaRawQm6WF(tSs6JTBnsDJvMaRawQm6WF), .Q7D2KKVRLkwEPktPhyCkSD(Q7D2KKVRLkwEPktPhyCkSD), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .OJ8T6Dl8xEKAEoVpEfestB(OJ8T6Dl8xEKAEoVpEfestB), .LsWvBUKOjIJIwF6hGU5kRC(LsWvBUKOjIJIwF6hGU5kRC) ); Ji2U3EhRqviNuqc0S23vUB AHBx0ZlFUu1jkAoPP4dmvG (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .OJ8T6Dl8xEKAEoVpEfestB(OJ8T6Dl8xEKAEoVpEfestB), .LsWvBUKOjIJIwF6hGU5kRC(LsWvBUKOjIJIwF6hGU5kRC), .QWAACQosHJOUrDgm1wJeoG(QWAACQosHJOUrDgm1wJeoG), .WgU2KCxd1j6m3EUCPiuf1F(WgU2KCxd1j6m3EUCPiuf1F), .y9Hu20tqKGzmg7O1xqeuAZH(y9Hu20tqKGzmg7O1xqeuAZH), .F9FfK0xrG2zVVJqYJzgfxD(F9FfK0xrG2zVVJqYJzgfxD), .xGMN0H1JXsbMHEVz1iuteB(xGMN0H1JXsbMHEVz1iuteB), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .E9kfQ0vBTIumIk9ATubhJH(E9kfQ0vBTIumIk9ATubhJH), .GFkF4uUefeRBOH9Wes3V5D(GFkF4uUefeRBOH9Wes3V5D) ); kFEYb0VSrycuLlb9yF6JYC O54bVOXwDTKIOcMLJdqYkE (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .NdNevEoWljk83nSbsGDU1C(NdNevEoWljk83nSbsGDU1C), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .Tf0EDmJTni9HuTSAYQFT2F(Tf0EDmJTni9HuTSAYQFT2F), .qp9pmnimi6dV0X7tI2Wt6B(qp9pmnimi6dV0X7tI2Wt6B) ); WTtof2St1Uu89F7e1eVXwF istKfX5aHEcknv2DxKn1PG (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .NdNevEoWljk83nSbsGDU1C(NdNevEoWljk83nSbsGDU1C), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .Gw5sPQAOzFLVF06eF1AOGF(Gw5sPQAOzFLVF06eF1AOGF), .uO7PvkjtbrbcoMU62rs5JF(uO7PvkjtbrbcoMU62rs5JF) ); bLNpla6dKRnNqV9xT7W46B WvEDazedW84qoYNTmNAHeB (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .S6Ue4SxCiz8dBHTO2guOUE(S6Ue4SxCiz8dBHTO2guOUE), .POhLmCr6emegQDte8TzyQ(POhLmCr6emegQDte8TzyQ), .E9kfQ0vBTIumIk9ATubhJH(E9kfQ0vBTIumIk9ATubhJH), .GFkF4uUefeRBOH9Wes3V5D(GFkF4uUefeRBOH9Wes3V5D), .NdNevEoWljk83nSbsGDU1C(NdNevEoWljk83nSbsGDU1C), .Tf0EDmJTni9HuTSAYQFT2F(Tf0EDmJTni9HuTSAYQFT2F), .qp9pmnimi6dV0X7tI2Wt6B(qp9pmnimi6dV0X7tI2Wt6B), .Gw5sPQAOzFLVF06eF1AOGF(Gw5sPQAOzFLVF06eF1AOGF), .uO7PvkjtbrbcoMU62rs5JF(uO7PvkjtbrbcoMU62rs5JF), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .qmhLAZZAHFrO09l1zXnPRC(qmhLAZZAHFrO09l1zXnPRC), .JMtgCMT5TVzyJSn9uILA1(JMtgCMT5TVzyJSn9uILA1), .xYJCS7zMCKI1yYR3Bx1XrD(xYJCS7zMCKI1yYR3Bx1XrD), .AaqUpSvCGAV1YR86nIsLWH(AaqUpSvCGAV1YR86nIsLWH) ); CcegpoX8iivyKlrAI1PDCD x21eZMV7RCoqI4FsDnz5jy (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .EnlAo7K66kKuzHIKWLmc1F(EnlAo7K66kKuzHIKWLmc1F), .ew3EeLap6s8rXmNrsqaTWH(ew3EeLap6s8rXmNrsqaTWH), .qmhLAZZAHFrO09l1zXnPRC(qmhLAZZAHFrO09l1zXnPRC), .JMtgCMT5TVzyJSn9uILA1(JMtgCMT5TVzyJSn9uILA1), .Z7ZDy0EvwvoCh1zahAqvSF(Z7ZDy0EvwvoCh1zahAqvSF), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .B58twvtfgVWGK5P29KavtH(B58twvtfgVWGK5P29KavtH), .qhk6Uhwhppvpssqm7Nh6XE(qhk6Uhwhppvpssqm7Nh6XE), .k3VfrgkD6DWITJL9WW5W4D(k3VfrgkD6DWITJL9WW5W4D), .pPn6MVGqBLqJ0xzN2WYfFG(pPn6MVGqBLqJ0xzN2WYfFG), .jNZ4xylBKAANfCL11XNxzB(jNZ4xylBKAANfCL11XNxzB) ); am04sFwquwsZE10aTKfoWG RpofGuiapIL2Va1hyZ1WGF (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .IPh1M0O3x0ioGlon72MROG(IPh1M0O3x0ioGlon72MROG), .Mt05SNCQbo0cCPNa1yEFyF(Mt05SNCQbo0cCPNa1yEFyF), .xYJCS7zMCKI1yYR3Bx1XrD(xYJCS7zMCKI1yYR3Bx1XrD), .AaqUpSvCGAV1YR86nIsLWH(AaqUpSvCGAV1YR86nIsLWH), .Z7ZDy0EvwvoCh1zahAqvSF(Z7ZDy0EvwvoCh1zahAqvSF), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .VWSiqDgxQN9a2J7zRy3p4E(VWSiqDgxQN9a2J7zRy3p4E), .LhqlKpPzANkuN2xC8HYciC(LhqlKpPzANkuN2xC8HYciC), .OUMqBzkN19EDa2VTABMa2E(OUMqBzkN19EDa2VTABMa2E), .qbEnMIxMUsx8pYkF1gFd7D(qbEnMIxMUsx8pYkF1gFd7D) ); ZW22u2kRuMcm5k35Olj0QH QMbS7KqGgbYlmDtgx5Wz1C (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .Ebx0yJLDGKevxkqzRPIfvG(Ebx0yJLDGKevxkqzRPIfvG), .B58twvtfgVWGK5P29KavtH(B58twvtfgVWGK5P29KavtH), .qhk6Uhwhppvpssqm7Nh6XE(qhk6Uhwhppvpssqm7Nh6XE), .VWSiqDgxQN9a2J7zRy3p4E(VWSiqDgxQN9a2J7zRy3p4E), .LhqlKpPzANkuN2xC8HYciC(LhqlKpPzANkuN2xC8HYciC), .jNZ4xylBKAANfCL11XNxzB(jNZ4xylBKAANfCL11XNxzB), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .A5SQIaNgqW7DcTqQkKRVeD(A5SQIaNgqW7DcTqQkKRVeD), .GaetbCaMty7UkzjqNoYErC(GaetbCaMty7UkzjqNoYErC), .k3VfrgkD6DWITJL9WW5W4D(M5AqS9R7rFTkWxwo8io2rH), .pPn6MVGqBLqJ0xzN2WYfFG(lcJo4MnEaj41ofRAtLkn4D), .iyuklaABkAlPLEQPPmVPCD(iyuklaABkAlPLEQPPmVPCD) ); assign mdal5obekPJm0ao7ZiZ4cF = A5SQIaNgqW7DcTqQkKRVeD; assign q4mhS1P9mOTwehAXXNmhxF = M5AqS9R7rFTkWxwo8io2rH; assign j8MMagsoA5t6IysA2ZD3X4F = 1'b1; u8mpVKkP8VQEVoiZ86piTAD bCLV4Qfl1BCm5WdQGQcoFC (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .j8MMagsoA5t6IysA2ZD3X4F(j8MMagsoA5t6IysA2ZD3X4F), .k3VfrgkD6DWITJL9WW5W4D(k3VfrgkD6DWITJL9WW5W4D), .pPn6MVGqBLqJ0xzN2WYfFG(pPn6MVGqBLqJ0xzN2WYfFG), .OUMqBzkN19EDa2VTABMa2E(OUMqBzkN19EDa2VTABMa2E), .qbEnMIxMUsx8pYkF1gFd7D(qbEnMIxMUsx8pYkF1gFd7D), .jNZ4xylBKAANfCL11XNxzB(jNZ4xylBKAANfCL11XNxzB), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .VWSiqDgxQN9a2J7zRy3p4E(aydyoHsGbz0wVGlm34qlsB), .LhqlKpPzANkuN2xC8HYciC(H0BpAwmwCivCDsbLQ5qvCC), .s1N0USypDrc4xyzxc4XEMr(s1N0USypDrc4xyzxc4XEMr), .sZ7bCwrhIAA80IOhzh695(sZ7bCwrhIAA80IOhzh695) ); assign vyWRmDyKy2RVVIdRBtzV5F = aydyoHsGbz0wVGlm34qlsB; assign SRoFC9yIIwEIUwYpoyy0QF = s1N0USypDrc4xyzxc4XEMr; assign wpHiLzmis5ns3l38MddOzE = GaetbCaMty7UkzjqNoYErC; assign j963sPBld8mpm71sqcvb8WF = lcJo4MnEaj41ofRAtLkn4D; assign Ic4vfYy6jnxaw8uXI98INH = H0BpAwmwCivCDsbLQ5qvCC; assign x2KkW4HKTQgVBmVskDu4RD = sZ7bCwrhIAA80IOhzh695; assign g1D8wSsV4Ksuy5G0qxKYMs = iyuklaABkAlPLEQPPmVPCD; endmodule