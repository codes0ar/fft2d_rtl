`timescale 1 ns / 1 ns module Jwp87To0uCqWGVPIwhN8ED (v04pHKxyc2sPW047bbyUgE, JAMOfrNHxGSYDF0urqkLN, Y7Nx2PyXNCTBUqlHxdhnVC, w9tDlZkclLF2jmOsqVKqWE, R6zf5iqRNVEGVBO8egq8kF, u5bboUjXYRZBbt1duYbKTG, mir92X5UlUGvLQSXmCuq9, hOMBB3qOa4Z6E9dukDYA0F); input v04pHKxyc2sPW047bbyUgE; input JAMOfrNHxGSYDF0urqkLN; input Y7Nx2PyXNCTBUqlHxdhnVC; input w9tDlZkclLF2jmOsqVKqWE; input R6zf5iqRNVEGVBO8egq8kF; output [6:0] u5bboUjXYRZBbt1duYbKTG; output mir92X5UlUGvLQSXmCuq9; output hOMBB3qOa4Z6E9dukDYA0F; reg [6:0] JomiEQo6ylRrlhLJPFsQTG; reg [1:0] X7FJ0jgk6hqdMN8BingGvE; reg [1:0] WXS42gmgDxS46057b3AGD; reg [6:0] GP01IUV0xObQQCSdqL463C; reg pDYTWTp6fyrEdA1XnDiP6E; reg [1:0] mb13NdjIe7rpJDLNih8AaE; reg Xf88wK4mkniJ6qfkmOXy2C; reg [6:0] i2IIQfdSjOGJ0HAlaZdYe; reg [1:0] xSW8arCNXsyV5zIEXuGUQB; reg [1:0] ck9Ya76HU61qWvvl3qwfRG; reg [6:0] dQhJtS5aSGZCPWaJqkkHi; reg t69iUVjqBKXZw2tNuE5YceG; reg [1:0] BNI9VucWF1TWsCAM4sBCHE; reg EIfu64RX7LMQGnynQeCGuD; reg [6:0] dsX1vjalwi3qczkXp6qk4; reg XMj0u82ecKWXG1WVNm9rRD; reg f72YcpkvfBqRpSxF9XKLJD; reg ZQj9wqlVlCJSDy0viA704C; wire B0yrqdBaR0HooAGUcvrwQB; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : h6oTzWU1a3otHwaiji95ID if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin JomiEQo6ylRrlhLJPFsQTG <= 7'b0000000; GP01IUV0xObQQCSdqL463C <= 7'b0000000; X7FJ0jgk6hqdMN8BingGvE <= 2'b00; WXS42gmgDxS46057b3AGD <= 2'b00; mb13NdjIe7rpJDLNih8AaE <= 2'b00; pDYTWTp6fyrEdA1XnDiP6E <= 1'b0; Xf88wK4mkniJ6qfkmOXy2C <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin JomiEQo6ylRrlhLJPFsQTG <= 7'b0000000; GP01IUV0xObQQCSdqL463C <= 7'b0000000; X7FJ0jgk6hqdMN8BingGvE <= 2'b00; WXS42gmgDxS46057b3AGD <= 2'b00; mb13NdjIe7rpJDLNih8AaE <= 2'b00; pDYTWTp6fyrEdA1XnDiP6E <= 1'b0; Xf88wK4mkniJ6qfkmOXy2C <= 1'b0; end else begin JomiEQo6ylRrlhLJPFsQTG <= i2IIQfdSjOGJ0HAlaZdYe; X7FJ0jgk6hqdMN8BingGvE <= xSW8arCNXsyV5zIEXuGUQB; WXS42gmgDxS46057b3AGD <= ck9Ya76HU61qWvvl3qwfRG; GP01IUV0xObQQCSdqL463C <= dQhJtS5aSGZCPWaJqkkHi; pDYTWTp6fyrEdA1XnDiP6E <= t69iUVjqBKXZw2tNuE5YceG; mb13NdjIe7rpJDLNih8AaE <= BNI9VucWF1TWsCAM4sBCHE; Xf88wK4mkniJ6qfkmOXy2C <= EIfu64RX7LMQGnynQeCGuD; end end end always @(GP01IUV0xObQQCSdqL463C, JomiEQo6ylRrlhLJPFsQTG, WXS42gmgDxS46057b3AGD, X7FJ0jgk6hqdMN8BingGvE, Xf88wK4mkniJ6qfkmOXy2C, Y7Nx2PyXNCTBUqlHxdhnVC, mb13NdjIe7rpJDLNih8AaE, pDYTWTp6fyrEdA1XnDiP6E, w9tDlZkclLF2jmOsqVKqWE) begin i2IIQfdSjOGJ0HAlaZdYe = JomiEQo6ylRrlhLJPFsQTG; xSW8arCNXsyV5zIEXuGUQB = X7FJ0jgk6hqdMN8BingGvE; ck9Ya76HU61qWvvl3qwfRG = WXS42gmgDxS46057b3AGD; dQhJtS5aSGZCPWaJqkkHi = GP01IUV0xObQQCSdqL463C; t69iUVjqBKXZw2tNuE5YceG = pDYTWTp6fyrEdA1XnDiP6E; BNI9VucWF1TWsCAM4sBCHE = mb13NdjIe7rpJDLNih8AaE; EIfu64RX7LMQGnynQeCGuD = Xf88wK4mkniJ6qfkmOXy2C; case ( mb13NdjIe7rpJDLNih8AaE) 2'b00 : begin BNI9VucWF1TWsCAM4sBCHE = 2'b00; EIfu64RX7LMQGnynQeCGuD = 1'b0; if (WXS42gmgDxS46057b3AGD == 2'b01) begin BNI9VucWF1TWsCAM4sBCHE = 2'b01; end end 2'b01 : begin EIfu64RX7LMQGnynQeCGuD = 1'b0; if (WXS42gmgDxS46057b3AGD == 2'b10) begin BNI9VucWF1TWsCAM4sBCHE = 2'b10; end end 2'b10 : begin EIfu64RX7LMQGnynQeCGuD = 1'b0; if (WXS42gmgDxS46057b3AGD == 2'b01) begin BNI9VucWF1TWsCAM4sBCHE = 2'b11; EIfu64RX7LMQGnynQeCGuD = 1'b1; end end 2'b11 : begin if (WXS42gmgDxS46057b3AGD == 2'b01) begin BNI9VucWF1TWsCAM4sBCHE = 2'b11; EIfu64RX7LMQGnynQeCGuD = 1'b1; end else begin EIfu64RX7LMQGnynQeCGuD = 1'b0; BNI9VucWF1TWsCAM4sBCHE = 2'b00; end end default : begin BNI9VucWF1TWsCAM4sBCHE = 2'b00; EIfu64RX7LMQGnynQeCGuD = 1'b0; end endcase case ( WXS42gmgDxS46057b3AGD) 2'b00 : begin ck9Ya76HU61qWvvl3qwfRG = 2'b00; dQhJtS5aSGZCPWaJqkkHi = 7'b0000000; XMj0u82ecKWXG1WVNm9rRD = 1'b0; if (Y7Nx2PyXNCTBUqlHxdhnVC && (JomiEQo6ylRrlhLJPFsQTG == 7'b1111111)) begin ck9Ya76HU61qWvvl3qwfRG = 2'b01; end end 2'b01 : begin ck9Ya76HU61qWvvl3qwfRG = 2'b01; XMj0u82ecKWXG1WVNm9rRD = w9tDlZkclLF2jmOsqVKqWE; if (w9tDlZkclLF2jmOsqVKqWE) begin if (GP01IUV0xObQQCSdqL463C == 7'b1111111) begin ck9Ya76HU61qWvvl3qwfRG = 2'b10; end dQhJtS5aSGZCPWaJqkkHi = GP01IUV0xObQQCSdqL463C + 7'b0000001; end end 2'b10 : begin XMj0u82ecKWXG1WVNm9rRD = 1'b1; if (GP01IUV0xObQQCSdqL463C == 7'b1111111) begin if (Y7Nx2PyXNCTBUqlHxdhnVC && (JomiEQo6ylRrlhLJPFsQTG == 7'b1111111)) begin ck9Ya76HU61qWvvl3qwfRG = 2'b01; end else begin ck9Ya76HU61qWvvl3qwfRG = 2'b00; end end dQhJtS5aSGZCPWaJqkkHi = GP01IUV0xObQQCSdqL463C + 7'b0000001; end default : begin ck9Ya76HU61qWvvl3qwfRG = 2'b00; dQhJtS5aSGZCPWaJqkkHi = 7'b0000000; XMj0u82ecKWXG1WVNm9rRD = 1'b0; end endcase case ( X7FJ0jgk6hqdMN8BingGvE) 2'b00 : begin xSW8arCNXsyV5zIEXuGUQB = 2'b00; i2IIQfdSjOGJ0HAlaZdYe = 7'b0000000; t69iUVjqBKXZw2tNuE5YceG = 1'b0; if (Y7Nx2PyXNCTBUqlHxdhnVC) begin xSW8arCNXsyV5zIEXuGUQB = 2'b01; i2IIQfdSjOGJ0HAlaZdYe = 7'b0000001; end end 2'b01 : begin xSW8arCNXsyV5zIEXuGUQB = 2'b01; t69iUVjqBKXZw2tNuE5YceG = 1'b0; if (Y7Nx2PyXNCTBUqlHxdhnVC) begin if (JomiEQo6ylRrlhLJPFsQTG == 7'b1111111) begin xSW8arCNXsyV5zIEXuGUQB = 2'b10; t69iUVjqBKXZw2tNuE5YceG = 1'b1; end else begin xSW8arCNXsyV5zIEXuGUQB = 2'b01; end i2IIQfdSjOGJ0HAlaZdYe = JomiEQo6ylRrlhLJPFsQTG + 7'b0000001; end end 2'b10 : begin xSW8arCNXsyV5zIEXuGUQB = 2'b10; if (Y7Nx2PyXNCTBUqlHxdhnVC) begin if (JomiEQo6ylRrlhLJPFsQTG == 7'b1111111) begin xSW8arCNXsyV5zIEXuGUQB = 2'b01; t69iUVjqBKXZw2tNuE5YceG = 1'b0; end else begin xSW8arCNXsyV5zIEXuGUQB = 2'b10; t69iUVjqBKXZw2tNuE5YceG = 1'b1; end i2IIQfdSjOGJ0HAlaZdYe = JomiEQo6ylRrlhLJPFsQTG + 7'b0000001; end end default : begin xSW8arCNXsyV5zIEXuGUQB = 2'b00; i2IIQfdSjOGJ0HAlaZdYe = 7'b1111111; t69iUVjqBKXZw2tNuE5YceG = 1'b0; end endcase dsX1vjalwi3qczkXp6qk4 = GP01IUV0xObQQCSdqL463C; f72YcpkvfBqRpSxF9XKLJD = pDYTWTp6fyrEdA1XnDiP6E; ZQj9wqlVlCJSDy0viA704C = Xf88wK4mkniJ6qfkmOXy2C; end assign u5bboUjXYRZBbt1duYbKTG = dsX1vjalwi3qczkXp6qk4; assign mir92X5UlUGvLQSXmCuq9 = XMj0u82ecKWXG1WVNm9rRD; assign hOMBB3qOa4Z6E9dukDYA0F = f72YcpkvfBqRpSxF9XKLJD; endmodule