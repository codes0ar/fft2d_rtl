`timescale 1 ns / 1 ns module IT7y3HrJPu7teNsd6CIHy (v04pHKxyc2sPW047bbyUgE, JAMOfrNHxGSYDF0urqkLN, OAkG388GVoqfAFfrsC3Z3, DP58bSOk4VSBFH6tnqlVTH, Ck459KQ1C8vRbine3lrkt, MCqIdNMOB0Mg1cefHLMjpH, j41GwwL8b9NI9l6ZScQ1PbG, i8H7HzN3cvjFks6MZ5qaqF, SAcShGLK2YZQrWHGqGVvjD, R6zf5iqRNVEGVBO8egq8kF, oEtRmwXRZkMV2JHZdumYM, ABAJKgUy1j1LH4rwhRtEnG); input v04pHKxyc2sPW047bbyUgE; input JAMOfrNHxGSYDF0urqkLN; input signed [15:0] OAkG388GVoqfAFfrsC3Z3; input signed [15:0] DP58bSOk4VSBFH6tnqlVTH; input Ck459KQ1C8vRbine3lrkt; input [1:0] MCqIdNMOB0Mg1cefHLMjpH; input j41GwwL8b9NI9l6ZScQ1PbG; input i8H7HzN3cvjFks6MZ5qaqF; input SAcShGLK2YZQrWHGqGVvjD; input R6zf5iqRNVEGVBO8egq8kF; output signed [15:0] oEtRmwXRZkMV2JHZdumYM; output signed [15:0] ABAJKgUy1j1LH4rwhRtEnG; wire UDLc9rLD6z9OmDzbHMGaFH; wire p34yBFVMhzZZL6P4BoBnpNE; wire yeU2ByaswMHNqD62x1WsFE; reg de21duRLbf27relCAO1YZB; reg cY321CCuBT3R7UOBs8HHRC; wire signed [15:0] iOhy3XYM3su7ndksftfCZG; wire [1:0] AECH0r3KnKo0RJFepDhYUD; wire twcuYIJzeZMBjyHmZ1FZDD; wire signed [15:0] dTkGd8OUQ83dmglc4Bt8vF; reg signed [15:0] d30z7znHID2VeOAFwdxJv3; wire signed [15:0] N2ZdE4zLlq5uRV4rcE2wdE; wire signed [15:0] csMK1iTp18g0vZYjmk9JZD; reg signed [15:0] BK42UUphOnOnQSjJxssa4C; reg YRZ5n25cqbkRRg7qQHehlC; reg FrWyM0cHsFwaFhwVURaveE; reg ONA2QGlNXG84z8xZQwVNBC; reg signed [16:0] peTrjdHrHks0XPmkydHeIE; reg signed [16:0] f5XQHcgrgY1gzEM7V5nLXsC; reg signed [16:0] h2pJbIsIwwtbYjPQ3REMsE; reg signed [16:0] m12eHWycKUWppJjZFhMLGB; reg signed [15:0] EBociv6W4lQ3ZvJNhw3Z8E; reg signed [15:0] TsaKCuYu0ALq2IfaWerghD; reg AZzMkYH85e704DYwHahVMC; reg signed [15:0] AOfQM5gh9zBuvl2vEIFejF; reg signed [15:0] c3emw2N1sQP4WZc39fVHCe; reg s2LfVOPizWwReFfjdJNWHmE; reg signed [15:0] D6SkVRQFbzIYRL1jZWDRY; reg signed [15:0] mbusDEwpxtjmRQrsdfHBrB; reg signed [15:0] a99DgeB7OWCpn91mJNssZhF; reg signed [15:0] h1qpvE4y6o27PpbIwHNDY0C; reg dPP1f4AA6YUsuLXPMqHOaD; reg g1C7IsBPLt2cJiWuoEetwG; reg GYoCMeSRAKsfSUDkd0UNSB; reg g6O7Lj8aAGN2KzWsHg2xoHG; reg signed [16:0] r9m0Z5zXiBEdpkbzXM3wtB; reg signed [16:0] FO3OGaIEzJ9wOWLjjp9nT; reg signed [16:0] NeoGTMM0QiM2bsdh1QoOLG; reg signed [16:0] XGDGyLQgR3aMe70DeSEyPG; reg signed [15:0] nREWllFEdkQ21QbMBOwhMF; reg signed [15:0] KKkNexVx5dAUwcjfJfUXrH; reg SYPfWJ9GCITBLgn5jpAhOB; reg signed [15:0] n3UlEbglw3m9cpZwISdPA5G; reg signed [15:0] tDiTrkLheWwDR0Ex16ijFG; reg LU1saL0hI4Ohy2cGQkKKG; reg signed [15:0] oPdwMlPCg2JbKLsFlPHvUF; reg signed [15:0] g4VHCMxNxJOHKs9dqZLxdG; reg signed [15:0] UMmIXixbRcgDTggJl4qF4C; reg signed [15:0] vLehpJq4NQsyWM0WolcfCF; reg w2dgPDpny5OW8JfhLyqq5VB; reg signed [15:0] mgknRxAcgFrHqTt5CZvnSF; reg signed [15:0] sCFM4WicR6deeSAdSwumP; reg BKNY6GzA6oGZumjzTATycD; reg signed [15:0] moYf2QENOIemSN5A51qCbG; reg signed [15:0] oLPVbqTEKvAQhOXQB7Fzp; reg ljAhzQENCBeBr4upZryUZB; reg signed [15:0] x9j7a5gok64zzNKnvdJNnE; reg signed [15:0] bPL0FcLvoxhO0amTUOV9QC; reg signed [15:0] r4JngA0ZVhEElGRZci9fohF; reg signed [15:0] a8xx20Fc5nKc8DbqSwNBuB; reg v9OrTxtIsmI18g6yKYT1kE; reg signed [16:0] kBrMhUdPuotKsdCeNoQ3DH; reg signed [16:0] G3Cb2SGcELdnfWn0LLaFIF; reg signed [16:0] HXNuTd4dJjyD0nq0PGZcbF; reg signed [16:0] Y2lV7uCKTIyXGwpwSv5xjF; reg signed [16:0] pckufEAGmvetxPhgoApe7D; reg signed [16:0] p9Op2WXQSnou9B2x2BL3j1B; reg signed [16:0] CeXlcosHh87Bq1wN4YYevD; reg signed [16:0] GI6VJV0Eq7K732wnimPfhF; reg signed [16:0] j9LCNq0jidDFu1rvmJmUKC; reg signed [16:0] k7Girg9LxT5XG1NL57rJ7hB; reg signed [16:0] q27eF7gVWuXwVP2KxqMHydB; reg signed [16:0] fQRY7P92irAHmLQDJuG00E; reg signed [16:0] N5IkIEUtQkHe2sBozuOXVE; reg signed [16:0] OPT67VtxcsDbilDQX22lNF; reg signed [16:0] uCz3oXsJUpbcNvG6iX2t9E; reg signed [16:0] m6EpxIuauHVhDE4hACkff9F; reg signed [16:0] fYwS5bgtgq2NnLZKEhMgS; reg signed [16:0] jrVFrTanH3gvKqaRhm37OD; reg signed [16:0] q0mjss3XEEQ5Du2vSLRk5CF; reg signed [16:0] s0qqNc1esXsOPKI0oAltk4; reg signed [16:0] RBQHsPk5GU0dXeqiTVc4lC; reg signed [16:0] CwJENrbhA04Cii9FbLO35; reg signed [16:0] IzmjnIjy7dTVYOBWEiIqXH; reg signed [16:0] kPYF09koGrRzabYjDQQY9F; reg signed [16:0] XMrIho4OvGjGyUn6NyRj2; reg signed [16:0] k0BAAYc1SrhTQTlkwXUFlhD; reg signed [16:0] ZaB7QLxBaJTFHQVpgVoZbH; reg signed [16:0] oD84amZL2f9PoEFtOiijQE; wire y47Mt5i1lVUvy3lpZgoyYhE; assign UDLc9rLD6z9OmDzbHMGaFH = Ck459KQ1C8vRbine3lrkt & i8H7HzN3cvjFks6MZ5qaqF; assign p34yBFVMhzZZL6P4BoBnpNE = ~ UDLc9rLD6z9OmDzbHMGaFH; assign yeU2ByaswMHNqD62x1WsFE = Ck459KQ1C8vRbine3lrkt & p34yBFVMhzZZL6P4BoBnpNE; always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : MczQYJ6MT1pYZD7C1UhQv if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin de21duRLbf27relCAO1YZB <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin de21duRLbf27relCAO1YZB <= 1'b0; end else begin de21duRLbf27relCAO1YZB <= j41GwwL8b9NI9l6ZScQ1PbG; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : xwyxj2YIc64Lxvl4r8S8mG if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin cY321CCuBT3R7UOBs8HHRC <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin cY321CCuBT3R7UOBs8HHRC <= 1'b0; end else begin cY321CCuBT3R7UOBs8HHRC <= de21duRLbf27relCAO1YZB; end end end PxGtD8RdpEuqNR1OqCny8D #(.AddrWidth(2), .DataWidth(16) ) BIK7TIfaOr4LLV21gmwOaE (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .E7QNJoK4KvAThVFhUlvl2G(iOhy3XYM3su7ndksftfCZG), .l30d1QakAt61ivcMw8sJQE(AECH0r3KnKo0RJFepDhYUD), .UKo8akspo4h0jsZ6g712NB(twcuYIJzeZMBjyHmZ1FZDD), .EYQG62ys4E6V8lISAdlW1C(MCqIdNMOB0Mg1cefHLMjpH), .HmVcl5yQin7hEovf3bwNG(dTkGd8OUQ83dmglc4Bt8vF) ); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : L1HBH8O5DRbGBa9XvBX70C if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin d30z7znHID2VeOAFwdxJv3 <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin d30z7znHID2VeOAFwdxJv3 <= 16'sb0000000000000000; end else begin d30z7znHID2VeOAFwdxJv3 <= dTkGd8OUQ83dmglc4Bt8vF; end end end PxGtD8RdpEuqNR1OqCny8D #(.AddrWidth(2), .DataWidth(16) ) y7YOcVduIzFPSAfkwovdwE (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .E7QNJoK4KvAThVFhUlvl2G(N2ZdE4zLlq5uRV4rcE2wdE), .l30d1QakAt61ivcMw8sJQE(AECH0r3KnKo0RJFepDhYUD), .UKo8akspo4h0jsZ6g712NB(twcuYIJzeZMBjyHmZ1FZDD), .EYQG62ys4E6V8lISAdlW1C(MCqIdNMOB0Mg1cefHLMjpH), .HmVcl5yQin7hEovf3bwNG(csMK1iTp18g0vZYjmk9JZD) ); always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : s2CWr6rrksK4W7N0omU97HD if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin BK42UUphOnOnQSjJxssa4C <= 16'sb0000000000000000; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin BK42UUphOnOnQSjJxssa4C <= 16'sb0000000000000000; end else begin BK42UUphOnOnQSjJxssa4C <= csMK1iTp18g0vZYjmk9JZD; end end end always @(posedge v04pHKxyc2sPW047bbyUgE or negedge JAMOfrNHxGSYDF0urqkLN) begin : xY29WdGpxj3QbNLuqj6PIH if (JAMOfrNHxGSYDF0urqkLN == 1'b0) begin YRZ5n25cqbkRRg7qQHehlC <= 1'b0; FrWyM0cHsFwaFhwVURaveE <= 1'b0; ONA2QGlNXG84z8xZQwVNBC <= 1'b0; peTrjdHrHks0XPmkydHeIE <= 17'sb00000000000000000; f5XQHcgrgY1gzEM7V5nLXsC <= 17'sb00000000000000000; h2pJbIsIwwtbYjPQ3REMsE <= 17'sb00000000000000000; m12eHWycKUWppJjZFhMLGB <= 17'sb00000000000000000; EBociv6W4lQ3ZvJNhw3Z8E <= 16'sb0000000000000000; TsaKCuYu0ALq2IfaWerghD <= 16'sb0000000000000000; AZzMkYH85e704DYwHahVMC <= 1'b0; AOfQM5gh9zBuvl2vEIFejF <= 16'sb0000000000000000; c3emw2N1sQP4WZc39fVHCe <= 16'sb0000000000000000; s2LfVOPizWwReFfjdJNWHmE <= 1'b0; D6SkVRQFbzIYRL1jZWDRY <= 16'sb0000000000000000; mbusDEwpxtjmRQrsdfHBrB <= 16'sb0000000000000000; a99DgeB7OWCpn91mJNssZhF <= 16'sb0000000000000000; h1qpvE4y6o27PpbIwHNDY0C <= 16'sb0000000000000000; dPP1f4AA6YUsuLXPMqHOaD <= 1'b0; end else begin if (R6zf5iqRNVEGVBO8egq8kF == 1'b1) begin YRZ5n25cqbkRRg7qQHehlC <= 1'b0; FrWyM0cHsFwaFhwVURaveE <= 1'b0; ONA2QGlNXG84z8xZQwVNBC <= 1'b0; peTrjdHrHks0XPmkydHeIE <= 17'sb00000000000000000; f5XQHcgrgY1gzEM7V5nLXsC <= 17'sb00000000000000000; h2pJbIsIwwtbYjPQ3REMsE <= 17'sb00000000000000000; m12eHWycKUWppJjZFhMLGB <= 17'sb00000000000000000; EBociv6W4lQ3ZvJNhw3Z8E <= 16'sb0000000000000000; TsaKCuYu0ALq2IfaWerghD <= 16'sb0000000000000000; AZzMkYH85e704DYwHahVMC <= 1'b0; AOfQM5gh9zBuvl2vEIFejF <= 16'sb0000000000000000; c3emw2N1sQP4WZc39fVHCe <= 16'sb0000000000000000; s2LfVOPizWwReFfjdJNWHmE <= 1'b0; D6SkVRQFbzIYRL1jZWDRY <= 16'sb0000000000000000; mbusDEwpxtjmRQrsdfHBrB <= 16'sb0000000000000000; a99DgeB7OWCpn91mJNssZhF <= 16'sb0000000000000000; h1qpvE4y6o27PpbIwHNDY0C <= 16'sb0000000000000000; dPP1f4AA6YUsuLXPMqHOaD <= 1'b0; end else begin YRZ5n25cqbkRRg7qQHehlC <= g1C7IsBPLt2cJiWuoEetwG; FrWyM0cHsFwaFhwVURaveE <= GYoCMeSRAKsfSUDkd0UNSB; ONA2QGlNXG84z8xZQwVNBC <= g6O7Lj8aAGN2KzWsHg2xoHG; peTrjdHrHks0XPmkydHeIE <= r9m0Z5zXiBEdpkbzXM3wtB; f5XQHcgrgY1gzEM7V5nLXsC <= FO3OGaIEzJ9wOWLjjp9nT; h2pJbIsIwwtbYjPQ3REMsE <= NeoGTMM0QiM2bsdh1QoOLG; m12eHWycKUWppJjZFhMLGB <= XGDGyLQgR3aMe70DeSEyPG; EBociv6W4lQ3ZvJNhw3Z8E <= nREWllFEdkQ21QbMBOwhMF; TsaKCuYu0ALq2IfaWerghD <= KKkNexVx5dAUwcjfJfUXrH; AZzMkYH85e704DYwHahVMC <= SYPfWJ9GCITBLgn5jpAhOB; AOfQM5gh9zBuvl2vEIFejF <= n3UlEbglw3m9cpZwISdPA5G; c3emw2N1sQP4WZc39fVHCe <= tDiTrkLheWwDR0Ex16ijFG; s2LfVOPizWwReFfjdJNWHmE <= LU1saL0hI4Ohy2cGQkKKG; D6SkVRQFbzIYRL1jZWDRY <= oPdwMlPCg2JbKLsFlPHvUF; mbusDEwpxtjmRQrsdfHBrB <= g4VHCMxNxJOHKs9dqZLxdG; a99DgeB7OWCpn91mJNssZhF <= UMmIXixbRcgDTggJl4qF4C; h1qpvE4y6o27PpbIwHNDY0C <= vLehpJq4NQsyWM0WolcfCF; dPP1f4AA6YUsuLXPMqHOaD <= w2dgPDpny5OW8JfhLyqq5VB; end end end always @(AOfQM5gh9zBuvl2vEIFejF, AZzMkYH85e704DYwHahVMC, BK42UUphOnOnQSjJxssa4C, D6SkVRQFbzIYRL1jZWDRY, DP58bSOk4VSBFH6tnqlVTH, EBociv6W4lQ3ZvJNhw3Z8E, FrWyM0cHsFwaFhwVURaveE, OAkG388GVoqfAFfrsC3Z3, ONA2QGlNXG84z8xZQwVNBC, SAcShGLK2YZQrWHGqGVvjD, TsaKCuYu0ALq2IfaWerghD, UDLc9rLD6z9OmDzbHMGaFH, YRZ5n25cqbkRRg7qQHehlC, a99DgeB7OWCpn91mJNssZhF, c3emw2N1sQP4WZc39fVHCe, cY321CCuBT3R7UOBs8HHRC, d30z7znHID2VeOAFwdxJv3, dPP1f4AA6YUsuLXPMqHOaD, f5XQHcgrgY1gzEM7V5nLXsC, h1qpvE4y6o27PpbIwHNDY0C, h2pJbIsIwwtbYjPQ3REMsE, m12eHWycKUWppJjZFhMLGB, mbusDEwpxtjmRQrsdfHBrB, peTrjdHrHks0XPmkydHeIE, s2LfVOPizWwReFfjdJNWHmE, yeU2ByaswMHNqD62x1WsFE) begin N5IkIEUtQkHe2sBozuOXVE = 17'sb00000000000000000; OPT67VtxcsDbilDQX22lNF = 17'sb00000000000000000; uCz3oXsJUpbcNvG6iX2t9E = 17'sb00000000000000000; m6EpxIuauHVhDE4hACkff9F = 17'sb00000000000000000; fYwS5bgtgq2NnLZKEhMgS = 17'sb00000000000000000; jrVFrTanH3gvKqaRhm37OD = 17'sb00000000000000000; q0mjss3XEEQ5Du2vSLRk5CF = 17'sb00000000000000000; s0qqNc1esXsOPKI0oAltk4 = 17'sb00000000000000000; RBQHsPk5GU0dXeqiTVc4lC = 17'sb00000000000000000; CwJENrbhA04Cii9FbLO35 = 17'sb00000000000000000; IzmjnIjy7dTVYOBWEiIqXH = 17'sb00000000000000000; kPYF09koGrRzabYjDQQY9F = 17'sb00000000000000000; XMrIho4OvGjGyUn6NyRj2 = 17'sb00000000000000000; k0BAAYc1SrhTQTlkwXUFlhD = 17'sb00000000000000000; ZaB7QLxBaJTFHQVpgVoZbH = 17'sb00000000000000000; oD84amZL2f9PoEFtOiijQE = 17'sb00000000000000000; r9m0Z5zXiBEdpkbzXM3wtB = peTrjdHrHks0XPmkydHeIE; FO3OGaIEzJ9wOWLjjp9nT = f5XQHcgrgY1gzEM7V5nLXsC; NeoGTMM0QiM2bsdh1QoOLG = h2pJbIsIwwtbYjPQ3REMsE; XGDGyLQgR3aMe70DeSEyPG = m12eHWycKUWppJjZFhMLGB; n3UlEbglw3m9cpZwISdPA5G = BK42UUphOnOnQSjJxssa4C; tDiTrkLheWwDR0Ex16ijFG = d30z7znHID2VeOAFwdxJv3; LU1saL0hI4Ohy2cGQkKKG = cY321CCuBT3R7UOBs8HHRC; nREWllFEdkQ21QbMBOwhMF = OAkG388GVoqfAFfrsC3Z3; KKkNexVx5dAUwcjfJfUXrH = DP58bSOk4VSBFH6tnqlVTH; SYPfWJ9GCITBLgn5jpAhOB = yeU2ByaswMHNqD62x1WsFE; g6O7Lj8aAGN2KzWsHg2xoHG = FrWyM0cHsFwaFhwVURaveE; GYoCMeSRAKsfSUDkd0UNSB = YRZ5n25cqbkRRg7qQHehlC; g1C7IsBPLt2cJiWuoEetwG = UDLc9rLD6z9OmDzbHMGaFH; if (dPP1f4AA6YUsuLXPMqHOaD) begin N5IkIEUtQkHe2sBozuOXVE = {BK42UUphOnOnQSjJxssa4C[15], BK42UUphOnOnQSjJxssa4C}; OPT67VtxcsDbilDQX22lNF = {h1qpvE4y6o27PpbIwHNDY0C[15], h1qpvE4y6o27PpbIwHNDY0C}; r9m0Z5zXiBEdpkbzXM3wtB = N5IkIEUtQkHe2sBozuOXVE + OPT67VtxcsDbilDQX22lNF; uCz3oXsJUpbcNvG6iX2t9E = {BK42UUphOnOnQSjJxssa4C[15], BK42UUphOnOnQSjJxssa4C}; m6EpxIuauHVhDE4hACkff9F = {h1qpvE4y6o27PpbIwHNDY0C[15], h1qpvE4y6o27PpbIwHNDY0C}; NeoGTMM0QiM2bsdh1QoOLG = uCz3oXsJUpbcNvG6iX2t9E - m6EpxIuauHVhDE4hACkff9F; fYwS5bgtgq2NnLZKEhMgS = {d30z7znHID2VeOAFwdxJv3[15], d30z7znHID2VeOAFwdxJv3}; jrVFrTanH3gvKqaRhm37OD = {a99DgeB7OWCpn91mJNssZhF[15], a99DgeB7OWCpn91mJNssZhF}; XGDGyLQgR3aMe70DeSEyPG = fYwS5bgtgq2NnLZKEhMgS + jrVFrTanH3gvKqaRhm37OD; q0mjss3XEEQ5Du2vSLRk5CF = {d30z7znHID2VeOAFwdxJv3[15], d30z7znHID2VeOAFwdxJv3}; s0qqNc1esXsOPKI0oAltk4 = {a99DgeB7OWCpn91mJNssZhF[15], a99DgeB7OWCpn91mJNssZhF}; FO3OGaIEzJ9wOWLjjp9nT = q0mjss3XEEQ5Du2vSLRk5CF - s0qqNc1esXsOPKI0oAltk4; end else begin RBQHsPk5GU0dXeqiTVc4lC = {BK42UUphOnOnQSjJxssa4C[15], BK42UUphOnOnQSjJxssa4C}; CwJENrbhA04Cii9FbLO35 = {a99DgeB7OWCpn91mJNssZhF[15], a99DgeB7OWCpn91mJNssZhF}; r9m0Z5zXiBEdpkbzXM3wtB = RBQHsPk5GU0dXeqiTVc4lC + CwJENrbhA04Cii9FbLO35; IzmjnIjy7dTVYOBWEiIqXH = {BK42UUphOnOnQSjJxssa4C[15], BK42UUphOnOnQSjJxssa4C}; kPYF09koGrRzabYjDQQY9F = {a99DgeB7OWCpn91mJNssZhF[15], a99DgeB7OWCpn91mJNssZhF}; NeoGTMM0QiM2bsdh1QoOLG = IzmjnIjy7dTVYOBWEiIqXH - kPYF09koGrRzabYjDQQY9F; XMrIho4OvGjGyUn6NyRj2 = {d30z7znHID2VeOAFwdxJv3[15], d30z7znHID2VeOAFwdxJv3}; k0BAAYc1SrhTQTlkwXUFlhD = {h1qpvE4y6o27PpbIwHNDY0C[15], h1qpvE4y6o27PpbIwHNDY0C}; FO3OGaIEzJ9wOWLjjp9nT = XMrIho4OvGjGyUn6NyRj2 + k0BAAYc1SrhTQTlkwXUFlhD; ZaB7QLxBaJTFHQVpgVoZbH = {d30z7znHID2VeOAFwdxJv3[15], d30z7znHID2VeOAFwdxJv3}; oD84amZL2f9PoEFtOiijQE = {h1qpvE4y6o27PpbIwHNDY0C[15], h1qpvE4y6o27PpbIwHNDY0C}; XGDGyLQgR3aMe70DeSEyPG = ZaB7QLxBaJTFHQVpgVoZbH - oD84amZL2f9PoEFtOiijQE; end UMmIXixbRcgDTggJl4qF4C = D6SkVRQFbzIYRL1jZWDRY; vLehpJq4NQsyWM0WolcfCF = mbusDEwpxtjmRQrsdfHBrB; oPdwMlPCg2JbKLsFlPHvUF = OAkG388GVoqfAFfrsC3Z3; g4VHCMxNxJOHKs9dqZLxdG = DP58bSOk4VSBFH6tnqlVTH; w2dgPDpny5OW8JfhLyqq5VB = SAcShGLK2YZQrWHGqGVvjD; mgknRxAcgFrHqTt5CZvnSF = AOfQM5gh9zBuvl2vEIFejF; sCFM4WicR6deeSAdSwumP = c3emw2N1sQP4WZc39fVHCe; BKNY6GzA6oGZumjzTATycD = s2LfVOPizWwReFfjdJNWHmE; moYf2QENOIemSN5A51qCbG = EBociv6W4lQ3ZvJNhw3Z8E; oLPVbqTEKvAQhOXQB7Fzp = TsaKCuYu0ALq2IfaWerghD; ljAhzQENCBeBr4upZryUZB = AZzMkYH85e704DYwHahVMC; kBrMhUdPuotKsdCeNoQ3DH = ({peTrjdHrHks0XPmkydHeIE[16], peTrjdHrHks0XPmkydHeIE[16:1]}) + $signed({1'b0, peTrjdHrHks0XPmkydHeIE[0]}); G3Cb2SGcELdnfWn0LLaFIF = kBrMhUdPuotKsdCeNoQ3DH >>> 8'd1; HXNuTd4dJjyD0nq0PGZcbF = {G3Cb2SGcELdnfWn0LLaFIF[15:0], 1'b0}; x9j7a5gok64zzNKnvdJNnE = HXNuTd4dJjyD0nq0PGZcbF[15:0]; Y2lV7uCKTIyXGwpwSv5xjF = ({f5XQHcgrgY1gzEM7V5nLXsC[16], f5XQHcgrgY1gzEM7V5nLXsC[16:1]}) + $signed({1'b0, f5XQHcgrgY1gzEM7V5nLXsC[0]}); pckufEAGmvetxPhgoApe7D = Y2lV7uCKTIyXGwpwSv5xjF >>> 8'd1; p9Op2WXQSnou9B2x2BL3j1B = {pckufEAGmvetxPhgoApe7D[15:0], 1'b0}; bPL0FcLvoxhO0amTUOV9QC = p9Op2WXQSnou9B2x2BL3j1B[15:0]; CeXlcosHh87Bq1wN4YYevD = ({h2pJbIsIwwtbYjPQ3REMsE[16], h2pJbIsIwwtbYjPQ3REMsE[16:1]}) + $signed({1'b0, h2pJbIsIwwtbYjPQ3REMsE[0]}); GI6VJV0Eq7K732wnimPfhF = CeXlcosHh87Bq1wN4YYevD >>> 8'd1; j9LCNq0jidDFu1rvmJmUKC = {GI6VJV0Eq7K732wnimPfhF[15:0], 1'b0}; r4JngA0ZVhEElGRZci9fohF = j9LCNq0jidDFu1rvmJmUKC[15:0]; k7Girg9LxT5XG1NL57rJ7hB = ({m12eHWycKUWppJjZFhMLGB[16], m12eHWycKUWppJjZFhMLGB[16:1]}) + $signed({1'b0, m12eHWycKUWppJjZFhMLGB[0]}); q27eF7gVWuXwVP2KxqMHydB = k7Girg9LxT5XG1NL57rJ7hB >>> 8'd1; fQRY7P92irAHmLQDJuG00E = {q27eF7gVWuXwVP2KxqMHydB[15:0], 1'b0}; a8xx20Fc5nKc8DbqSwNBuB = fQRY7P92irAHmLQDJuG00E[15:0]; v9OrTxtIsmI18g6yKYT1kE = ONA2QGlNXG84z8xZQwVNBC; end CF9h42pdrNtczTiNIr4DCB VmvCiKePrWgzRko4o2171 (.v04pHKxyc2sPW047bbyUgE(v04pHKxyc2sPW047bbyUgE), .JAMOfrNHxGSYDF0urqkLN(JAMOfrNHxGSYDF0urqkLN), .Ck459KQ1C8vRbine3lrkt(Ck459KQ1C8vRbine3lrkt), .mgknRxAcgFrHqTt5CZvnSF(mgknRxAcgFrHqTt5CZvnSF), .sCFM4WicR6deeSAdSwumP(sCFM4WicR6deeSAdSwumP), .BKNY6GzA6oGZumjzTATycD(BKNY6GzA6oGZumjzTATycD), .moYf2QENOIemSN5A51qCbG(moYf2QENOIemSN5A51qCbG), .oLPVbqTEKvAQhOXQB7Fzp(oLPVbqTEKvAQhOXQB7Fzp), .ljAhzQENCBeBr4upZryUZB(ljAhzQENCBeBr4upZryUZB), .x9j7a5gok64zzNKnvdJNnE(x9j7a5gok64zzNKnvdJNnE), .bPL0FcLvoxhO0amTUOV9QC(bPL0FcLvoxhO0amTUOV9QC), .r4JngA0ZVhEElGRZci9fohF(r4JngA0ZVhEElGRZci9fohF), .a8xx20Fc5nKc8DbqSwNBuB(a8xx20Fc5nKc8DbqSwNBuB), .v9OrTxtIsmI18g6yKYT1kE(v9OrTxtIsmI18g6yKYT1kE), .R6zf5iqRNVEGVBO8egq8kF(R6zf5iqRNVEGVBO8egq8kF), .N2ZdE4zLlq5uRV4rcE2wdE(N2ZdE4zLlq5uRV4rcE2wdE), .iOhy3XYM3su7ndksftfCZG(iOhy3XYM3su7ndksftfCZG), .AECH0r3KnKo0RJFepDhYUD(AECH0r3KnKo0RJFepDhYUD), .twcuYIJzeZMBjyHmZ1FZDD(twcuYIJzeZMBjyHmZ1FZDD), .oEtRmwXRZkMV2JHZdumYM(oEtRmwXRZkMV2JHZdumYM), .ABAJKgUy1j1LH4rwhRtEnG(ABAJKgUy1j1LH4rwhRtEnG) ); endmodule