`timescale 1 ns / 1 ns module e8HeF7GSPxfrhisMVdBBvN (yQNwAzareGOhTeFAcGgFWE, jqBlsvEQIekR8Gt2pzz5n); input [31:0] yQNwAzareGOhTeFAcGgFWE; output [15:0] jqBlsvEQIekR8Gt2pzz5n; wire [15:0] sBKdfayBUR3Ntuy7EQrBgD; wire [15:0] mOhSSytk7nWnNPtZQ4VYl; wire [15:0] Qs9FrBdvqkfYe6HDuZ5x4G; wire [15:0] KeIx4znJ7NwHTA7mczkoe; wire [15:0] pdFb2Ar1wmoFWvU07SJWFF; wire [15:0] QPMLNVTOMA3OrhKJ2KbGiH; wire [15:0] DFkPjhhRCMOYOsSbu6aQEF; wire [15:0] NtHjaHzNt0xelhyuxLFDIE; wire [15:0] vYbET88zhkForoawWcw18E; wire [15:0] x1hHF4Y8ZceMfdfnAWH8Mc; wire [15:0] Euq2kmsb9LTNk8IgXS0ol; wire [15:0] s3eHG7L1MH98LfVKO4py88F; wire [15:0] JBmdc6zOYDzlxqcx1YjZb; wire [15:0] zawXB1WtJmMfC1cNcABaaE; wire [15:0] nORSkpKN0CGUenzeTFfUDB; wire fXtzdo4P9yi1Ciqp6QBfjC; wire [15:0] ajv4lpvFjoE3ofDGMFu5cE; wire [15:0] fatWyfdkxQ7BzaNjbRT4QD; wire n7hoWcccdXrFN0C874HrpEB; wire [1:0] ebKSCnB4aCunFgmKuqoZYH; wire [15:0] GySsTihj2cPCBENEuIyCSD; wire [15:0] xkbuOVpB2WYtI1blvBLI4F; wire K3vG6BZkHRRw0KY26D9MZB; wire [1:0] lUScGnUZMrmRi9dRMz0LkD; wire [15:0] SrrYc2LpbOfxe2q5vcN0ZB; wire [15:0] HXKQBF1mrJNaqSvHX0NNjE; wire n9yUlIfpQp88T4XdCnh7CDF; wire [1:0] d5CXluM5YmRNluM6LdzEuRD; wire [15:0] NEJXc3NqgfPBnBXZhsnaBH; wire [15:0] pfAEfAzOvu7FtEVFulxbzD; wire JlM61doAjTFQp2IhAs1cSH; wire [1:0] gBkF6hCOJWWy5LuZbB48v; wire [15:0] Ndwbn1qn70dbIKd1eeGFLH; wire [15:0] w5i8Ug2h8McUnQb3WOIwnOC; wire yyuLRu89eNc5LwJryJc7rE; wire [1:0] gjjq7XRjRpkPoRKYu5l6n; wire [15:0] A4JsqN6vYZ3AEKxV7Ife2D; wire [15:0] jqLr7Qvd3gtCcUpcnS2jjE; wire ScrD9UeAxKjITzyoNx94zC; wire [1:0] ATVtgjciSvCRUI7H3Y9tuD; wire [15:0] kPPlhFE2ldEEQzJYYPeCpC; wire [15:0] f1vtztaLG8k7ETvXjGQi2D; wire WM76Z8aHuuoFAdf9WffSUE; wire [1:0] FBdqgz94a8SGX1FULhpnhF; wire [15:0] eq6ExCvRAypD8ZXX1hJg2G; wire [15:0] zqoHGtfy6Sfo7Yl3f754XE; wire TkIpU7Kfy1Dc33ZRJQj19C; wire [1:0] NtsaMyVZXVYmztcjOvOk8; wire [15:0] e1s8qm2TAAcsGxoTmde7BD; wire [15:0] PhcezgX6tOzisplfkIJwjD; wire a99cv4QPwIifb55QksH05aG; wire [1:0] q26YIydocFfUg15Xj6RX5F; wire [15:0] N3LfeWGStZMqNRoOruJiLB; wire [15:0] Rzd2KleDteHJnQGGQBspBG; wire rvf3v0TbKi0SUQyjoMm0WE; wire [1:0] K2KmCTF5G7ost89y9oqLiD; wire [15:0] c1ronCM2H01cjuP1wRFxc7C; wire [15:0] ue4zD618Z3SRCgWU1P9vMG; wire M9E8thmcmP8jFioTvkEhuB; wire [1:0] iUgDeFg7wK7VmcsUejECJE; wire [15:0] TKuu61vVE7qT0QqU65DVCB; wire [15:0] h75JuQ3GzF4Eyf7QEyVL2ND; wire taujhy7mQH8DNG1xOnzviE; wire [1:0] CzuyViL53TclNSqIDzrvkF; wire [15:0] UXVpiMug8SwGCNbjOrLnFH; wire [15:0] AdUKfM0WY49g0VXTwB2VgF; wire fqh7z20DXcDCXlGSq1hmlH; assign sBKdfayBUR3Ntuy7EQrBgD = yQNwAzareGOhTeFAcGgFWE[15:0]; assign mOhSSytk7nWnNPtZQ4VYl = 16'b0001000000000000; assign Qs9FrBdvqkfYe6HDuZ5x4G = 16'b0000100000000000; assign KeIx4znJ7NwHTA7mczkoe = 16'b0000010000000000; assign pdFb2Ar1wmoFWvU07SJWFF = 16'b0000001000000000; assign QPMLNVTOMA3OrhKJ2KbGiH = 16'b0000000100000000; assign DFkPjhhRCMOYOsSbu6aQEF = 16'b0000000010000000; assign NtHjaHzNt0xelhyuxLFDIE = 16'b0000000001000000; assign vYbET88zhkForoawWcw18E = 16'b0000000000100000; assign x1hHF4Y8ZceMfdfnAWH8Mc = 16'b0000000000010000; assign Euq2kmsb9LTNk8IgXS0ol = 16'b0000000000001000; assign s3eHG7L1MH98LfVKO4py88F = 16'b0000000000000100; assign JBmdc6zOYDzlxqcx1YjZb = 16'b0000000000000010; assign zawXB1WtJmMfC1cNcABaaE = 16'b0000000000000001; assign nORSkpKN0CGUenzeTFfUDB = sBKdfayBUR3Ntuy7EQrBgD & mOhSSytk7nWnNPtZQ4VYl; assign fXtzdo4P9yi1Ciqp6QBfjC = (|nORSkpKN0CGUenzeTFfUDB[15:0]); assign ajv4lpvFjoE3ofDGMFu5cE = {15'b0, fXtzdo4P9yi1Ciqp6QBfjC}; assign fatWyfdkxQ7BzaNjbRT4QD = sBKdfayBUR3Ntuy7EQrBgD & Qs9FrBdvqkfYe6HDuZ5x4G; assign n7hoWcccdXrFN0C874HrpEB = (|fatWyfdkxQ7BzaNjbRT4QD[15:0]); assign ebKSCnB4aCunFgmKuqoZYH = {1'b0, n7hoWcccdXrFN0C874HrpEB}; assign GySsTihj2cPCBENEuIyCSD = {13'b0, {ebKSCnB4aCunFgmKuqoZYH, 1'b0}}; assign xkbuOVpB2WYtI1blvBLI4F = sBKdfayBUR3Ntuy7EQrBgD & KeIx4znJ7NwHTA7mczkoe; assign K3vG6BZkHRRw0KY26D9MZB = (|xkbuOVpB2WYtI1blvBLI4F[15:0]); assign lUScGnUZMrmRi9dRMz0LkD = {1'b0, K3vG6BZkHRRw0KY26D9MZB}; assign SrrYc2LpbOfxe2q5vcN0ZB = {12'b0, {lUScGnUZMrmRi9dRMz0LkD, 2'b00}}; assign HXKQBF1mrJNaqSvHX0NNjE = sBKdfayBUR3Ntuy7EQrBgD & pdFb2Ar1wmoFWvU07SJWFF; assign n9yUlIfpQp88T4XdCnh7CDF = (|HXKQBF1mrJNaqSvHX0NNjE[15:0]); assign d5CXluM5YmRNluM6LdzEuRD = {1'b0, n9yUlIfpQp88T4XdCnh7CDF}; assign NEJXc3NqgfPBnBXZhsnaBH = {11'b0, {d5CXluM5YmRNluM6LdzEuRD, 3'b000}}; assign pfAEfAzOvu7FtEVFulxbzD = sBKdfayBUR3Ntuy7EQrBgD & QPMLNVTOMA3OrhKJ2KbGiH; assign JlM61doAjTFQp2IhAs1cSH = (|pfAEfAzOvu7FtEVFulxbzD[15:0]); assign gBkF6hCOJWWy5LuZbB48v = {1'b0, JlM61doAjTFQp2IhAs1cSH}; assign Ndwbn1qn70dbIKd1eeGFLH = {10'b0, {gBkF6hCOJWWy5LuZbB48v, 4'b0000}}; assign w5i8Ug2h8McUnQb3WOIwnOC = sBKdfayBUR3Ntuy7EQrBgD & DFkPjhhRCMOYOsSbu6aQEF; assign yyuLRu89eNc5LwJryJc7rE = (|w5i8Ug2h8McUnQb3WOIwnOC[15:0]); assign gjjq7XRjRpkPoRKYu5l6n = {1'b0, yyuLRu89eNc5LwJryJc7rE}; assign A4JsqN6vYZ3AEKxV7Ife2D = {9'b0, {gjjq7XRjRpkPoRKYu5l6n, 5'b00000}}; assign jqLr7Qvd3gtCcUpcnS2jjE = sBKdfayBUR3Ntuy7EQrBgD & NtHjaHzNt0xelhyuxLFDIE; assign ScrD9UeAxKjITzyoNx94zC = (|jqLr7Qvd3gtCcUpcnS2jjE[15:0]); assign ATVtgjciSvCRUI7H3Y9tuD = {1'b0, ScrD9UeAxKjITzyoNx94zC}; assign kPPlhFE2ldEEQzJYYPeCpC = {8'b0, {ATVtgjciSvCRUI7H3Y9tuD, 6'b000000}}; assign f1vtztaLG8k7ETvXjGQi2D = sBKdfayBUR3Ntuy7EQrBgD & vYbET88zhkForoawWcw18E; assign WM76Z8aHuuoFAdf9WffSUE = (|f1vtztaLG8k7ETvXjGQi2D[15:0]); assign FBdqgz94a8SGX1FULhpnhF = {1'b0, WM76Z8aHuuoFAdf9WffSUE}; assign eq6ExCvRAypD8ZXX1hJg2G = {7'b0, {FBdqgz94a8SGX1FULhpnhF, 7'b0000000}}; assign zqoHGtfy6Sfo7Yl3f754XE = sBKdfayBUR3Ntuy7EQrBgD & x1hHF4Y8ZceMfdfnAWH8Mc; assign TkIpU7Kfy1Dc33ZRJQj19C = (|zqoHGtfy6Sfo7Yl3f754XE[15:0]); assign NtsaMyVZXVYmztcjOvOk8 = {1'b0, TkIpU7Kfy1Dc33ZRJQj19C}; assign e1s8qm2TAAcsGxoTmde7BD = {6'b0, {NtsaMyVZXVYmztcjOvOk8, 8'b00000000}}; assign PhcezgX6tOzisplfkIJwjD = sBKdfayBUR3Ntuy7EQrBgD & Euq2kmsb9LTNk8IgXS0ol; assign a99cv4QPwIifb55QksH05aG = (|PhcezgX6tOzisplfkIJwjD[15:0]); assign q26YIydocFfUg15Xj6RX5F = {1'b0, a99cv4QPwIifb55QksH05aG}; assign N3LfeWGStZMqNRoOruJiLB = {5'b0, {q26YIydocFfUg15Xj6RX5F, 9'b000000000}}; assign Rzd2KleDteHJnQGGQBspBG = sBKdfayBUR3Ntuy7EQrBgD & s3eHG7L1MH98LfVKO4py88F; assign rvf3v0TbKi0SUQyjoMm0WE = (|Rzd2KleDteHJnQGGQBspBG[15:0]); assign K2KmCTF5G7ost89y9oqLiD = {1'b0, rvf3v0TbKi0SUQyjoMm0WE}; assign c1ronCM2H01cjuP1wRFxc7C = {4'b0, {K2KmCTF5G7ost89y9oqLiD, 10'b0000000000}}; assign ue4zD618Z3SRCgWU1P9vMG = sBKdfayBUR3Ntuy7EQrBgD & JBmdc6zOYDzlxqcx1YjZb; assign M9E8thmcmP8jFioTvkEhuB = (|ue4zD618Z3SRCgWU1P9vMG[15:0]); assign iUgDeFg7wK7VmcsUejECJE = {1'b0, M9E8thmcmP8jFioTvkEhuB}; assign TKuu61vVE7qT0QqU65DVCB = {3'b0, {iUgDeFg7wK7VmcsUejECJE, 11'b00000000000}}; assign h75JuQ3GzF4Eyf7QEyVL2ND = sBKdfayBUR3Ntuy7EQrBgD & zawXB1WtJmMfC1cNcABaaE; assign taujhy7mQH8DNG1xOnzviE = (|h75JuQ3GzF4Eyf7QEyVL2ND[15:0]); assign CzuyViL53TclNSqIDzrvkF = {1'b0, taujhy7mQH8DNG1xOnzviE}; assign UXVpiMug8SwGCNbjOrLnFH = {2'b0, {CzuyViL53TclNSqIDzrvkF, 12'b000000000000}}; assign AdUKfM0WY49g0VXTwB2VgF = UXVpiMug8SwGCNbjOrLnFH | (TKuu61vVE7qT0QqU65DVCB | (c1ronCM2H01cjuP1wRFxc7C | (N3LfeWGStZMqNRoOruJiLB | (e1s8qm2TAAcsGxoTmde7BD | (eq6ExCvRAypD8ZXX1hJg2G | (kPPlhFE2ldEEQzJYYPeCpC | (A4JsqN6vYZ3AEKxV7Ife2D | (Ndwbn1qn70dbIKd1eeGFLH | (NEJXc3NqgfPBnBXZhsnaBH | (SrrYc2LpbOfxe2q5vcN0ZB | (ajv4lpvFjoE3ofDGMFu5cE | GySsTihj2cPCBENEuIyCSD))))))))))); assign jqBlsvEQIekR8Gt2pzz5n = AdUKfM0WY49g0VXTwB2VgF; endmodule